library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- This contains 0.72 of the ICE T65 (a.k.a AtomCpuMon) firmware

-- For f_log2 definition
use WORK.SynthCtrlPack.all;

entity XPM is
    generic (
        WIDTH : integer;
        SIZE  : integer
    );
    port(
        cp2     : in  std_logic;
        ce      : in  std_logic;
        address : in  std_logic_vector(f_log2(SIZE) - 1 downto 0);
        din     : in  std_logic_vector(WIDTH - 1 downto 0);
        dout    : out std_logic_vector(WIDTH - 1 downto 0);
        we      : in  std_logic
    );
end;

architecture RTL of XPM is

    type ram_type is array (0 to SIZE - 1) of std_logic_vector (WIDTH - 1 downto 0);

    signal RAM : ram_type := (
        x"940C",
        x"042C",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"940C",
        x"044E",
        x"14B1",
        x"14B4",
        x"1578",
        x"14C3",
        x"14CF",
        x"14E3",
        x"14E8",
        x"14ED",
        x"14F7",
        x"14FC",
        x"14F2",
        x"1578",
        x"1501",
        x"1519",
        x"1531",
        x"1549",
        x"1561",
        x"6463",
        x"6E69",
        x"706F",
        x"7573",
        x"5878",
        x"005B",
        x"6E55",
        x"6E6B",
        x"776F",
        x"206E",
        x"6F63",
        x"6D6D",
        x"6E61",
        x"2064",
        x"7325",
        x"000A",
        x"6E49",
        x"6574",
        x"7272",
        x"7075",
        x"6574",
        x"0A64",
        x"4300",
        x"5550",
        x"6620",
        x"6572",
        x"2065",
        x"7572",
        x"6E6E",
        x"6E69",
        x"2E67",
        x"2E2E",
        x"000A",
        x"2020",
        x"2020",
        x"5825",
        x"3D20",
        x"2520",
        x"0A73",
        x"5400",
        x"6972",
        x"6767",
        x"7265",
        x"4320",
        x"646F",
        x"7365",
        x"0A3A",
        x"2000",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"5200",
        x"6D65",
        x"766F",
        x"6E69",
        x"2067",
        x"4E00",
        x"206F",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"6573",
        x"0A74",
        x"2900",
        x"000A",
        x"2820",
        x"2500",
        x"3A64",
        x"2520",
        x"3430",
        x"2058",
        x"616D",
        x"6B73",
        x"2520",
        x"3430",
        x"3A58",
        x"0020",
        x"6520",
        x"616E",
        x"6C62",
        x"6465",
        x"000A",
        x"6920",
        x"686E",
        x"6269",
        x"7469",
        x"6465",
        x"000A",
        x"7325",
        x"7300",
        x"696B",
        x"7070",
        x"6E69",
        x"2067",
        x"2553",
        x"0A64",
        x"7400",
        x"6172",
        x"736E",
        x"6566",
        x"7272",
        x"6465",
        x"2520",
        x"2064",
        x"7962",
        x"6574",
        x"2073",
        x"6F74",
        x"3020",
        x"2578",
        x"3430",
        x"2078",
        x"202D",
        x"7830",
        x"3025",
        x"7834",
        x"000A",
        x"6572",
        x"6963",
        x"7665",
        x"6465",
        x"2520",
        x"2064",
        x"6F67",
        x"646F",
        x"7220",
        x"6365",
        x"726F",
        x"7364",
        x"202C",
        x"6425",
        x"6220",
        x"6461",
        x"7220",
        x"6365",
        x"726F",
        x"7364",
        x"000A",
        x"6553",
        x"646E",
        x"6620",
        x"6C69",
        x"2065",
        x"6F6E",
        x"2E77",
        x"2E2E",
        x"000A",
        x"7263",
        x"3A63",
        x"2520",
        x"3430",
        x"0A58",
        x"5700",
        x"3A72",
        x"2520",
        x"3430",
        x"2058",
        x"6F74",
        x"2520",
        x"3430",
        x"2058",
        x"203D",
        x"3025",
        x"5832",
        x"000A",
        x"6E49",
        x"6574",
        x"7272",
        x"7075",
        x"6574",
        x"2064",
        x"6661",
        x"6574",
        x"2072",
        x"6C25",
        x"2064",
        x"6E69",
        x"7473",
        x"7572",
        x"7463",
        x"6F69",
        x"736E",
        x"000A",
        x"7453",
        x"7065",
        x"6970",
        x"676E",
        x"2520",
        x"646C",
        x"6920",
        x"736E",
        x"7274",
        x"6375",
        x"6974",
        x"6E6F",
        x"0A73",
        x"4E00",
        x"6D75",
        x"6562",
        x"2072",
        x"666F",
        x"6920",
        x"736E",
        x"7574",
        x"7463",
        x"6F69",
        x"736E",
        x"6D20",
        x"7375",
        x"2074",
        x"6562",
        x"7020",
        x"736F",
        x"7469",
        x"7669",
        x"0A65",
        x"2000",
        x"2020",
        x"2520",
        x"0A73",
        x"4300",
        x"6D6F",
        x"616D",
        x"646E",
        x"3A73",
        x"000A",
        x"6552",
        x"6573",
        x"7474",
        x"6E69",
        x"2067",
        x"5043",
        x"0A55",
        x"3A00",
        x"7020",
        x"7361",
        x"6573",
        x"0A64",
        x"3A00",
        x"6620",
        x"6961",
        x"656C",
        x"3A64",
        x"2520",
        x"2064",
        x"7265",
        x"6F72",
        x"7372",
        x"000A",
        x"2520",
        x"3230",
        x"0058",
        x"654D",
        x"6F6D",
        x"7972",
        x"7420",
        x"7365",
        x"3A74",
        x"2520",
        x"0073",
        x"6146",
        x"6C69",
        x"6120",
        x"2074",
        x"3025",
        x"6C34",
        x"2058",
        x"5728",
        x"6F72",
        x"6574",
        x"203A",
        x"3025",
        x"5832",
        x"202C",
        x"6552",
        x"6461",
        x"6220",
        x"6361",
        x"206B",
        x"3025",
        x"5832",
        x"0A29",
        x"2000",
        x"6C61",
        x"6572",
        x"6461",
        x"2079",
        x"6573",
        x"2074",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"4100",
        x"6C6C",
        x"2520",
        x"2064",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"7261",
        x"2065",
        x"6C61",
        x"6572",
        x"6461",
        x"2079",
        x"6573",
        x"0A74",
        x"2000",
        x"6573",
        x"2074",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"5400",
        x"6172",
        x"6963",
        x"676E",
        x"6420",
        x"7369",
        x"6261",
        x"656C",
        x"0A64",
        x"5400",
        x"6172",
        x"6963",
        x"676E",
        x"6520",
        x"6576",
        x"7972",
        x"2520",
        x"646C",
        x"6920",
        x"736E",
        x"7274",
        x"6375",
        x"6974",
        x"6E6F",
        x"2073",
        x"6877",
        x"6C69",
        x"2065",
        x"6973",
        x"676E",
        x"656C",
        x"7320",
        x"6574",
        x"7070",
        x"6E69",
        x"0A67",
        x"4200",
        x"6572",
        x"6B61",
        x"6F70",
        x"6E69",
        x"2F74",
        x"6177",
        x"6374",
        x"2068",
        x"6F6E",
        x"2074",
        x"6573",
        x"2074",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"2500",
        x"2064",
        x"6177",
        x"6374",
        x"6568",
        x"2F73",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"6D69",
        x"6C70",
        x"6D65",
        x"6E65",
        x"6574",
        x"0A64",
        x"4300",
        x"6D6F",
        x"6970",
        x"656C",
        x"2064",
        x"7461",
        x"2520",
        x"2073",
        x"6E6F",
        x"2520",
        x"0A73",
        x"2500",
        x"2073",
        x"6E49",
        x"432D",
        x"7269",
        x"7563",
        x"7469",
        x"4520",
        x"756D",
        x"616C",
        x"6F74",
        x"2072",
        x"6576",
        x"7372",
        x"6F69",
        x"206E",
        x"7325",
        x"000A",
        x"000A",
        x"7220",
        x"6165",
        x"6964",
        x"676E",
        x"2000",
        x"7277",
        x"7469",
        x"6E69",
        x"0067",
        x"6820",
        x"7469",
        x"6120",
        x"2074",
        x"3025",
        x"5834",
        x"7400",
        x"6972",
        x"6767",
        x"7265",
        x"203A",
        x"4C49",
        x"454C",
        x"4147",
        x"004C",
        x"7274",
        x"6769",
        x"6567",
        x"3A72",
        x"2520",
        x"0073",
        x"7325",
        x"2C00",
        x"0020",
        x"3025",
        x"6C32",
        x"2E64",
        x"3025",
        x"6C36",
        x"3A64",
        x"0020",
        x"6E49",
        x"6F63",
        x"736E",
        x"7369",
        x"6574",
        x"746E",
        x"5220",
        x"3A64",
        x"2520",
        x"3230",
        x"2058",
        x"3E3C",
        x"2520",
        x"3230",
        x"0A58",
        x"0A00",
        x"5200",
        x"3A64",
        x"0020",
        x"000A",
        x"7257",
        x"203A",
        x"0A00",
        x"2000",
        x"2500",
        x"3230",
        x"2058",
        x"2500",
        x"3430",
        x"2058",
        x"2000",
        x"3025",
        x"5834",
        x"3D20",
        x"2520",
        x"3230",
        x"2058",
        x"0020",
        x"6325",
        x"3E00",
        x"203E",
        x"1B00",
        x"305B",
        x"303B",
        x"0048",
        x"5B1B",
        x"4A32",
        x"1B00",
        x"305B",
        x"303B",
        x"0048",
        x"5B1B",
        x"4A32",
        x"0A00",
        x"2800",
        x"3025",
        x"5832",
        x"3025",
        x"5832",
        x"582C",
        x"0029",
        x"2528",
        x"3230",
        x"2558",
        x"3230",
        x"2958",
        x"2020",
        x"2500",
        x"3230",
        x"2558",
        x"3230",
        x"2C58",
        x"2059",
        x"0020",
        x"3025",
        x"5832",
        x"3025",
        x"5832",
        x"582C",
        x"2020",
        x"2500",
        x"3230",
        x"2558",
        x"3230",
        x"2058",
        x"2020",
        x"0020",
        x"2528",
        x"3230",
        x"2958",
        x"592C",
        x"2020",
        x"2800",
        x"3025",
        x"5832",
        x"582C",
        x"2029",
        x"0020",
        x"2528",
        x"3230",
        x"2958",
        x"2020",
        x"2020",
        x"2500",
        x"3230",
        x"2C58",
        x"2059",
        x"2020",
        x"0020",
        x"3025",
        x"5832",
        x"582C",
        x"2020",
        x"2020",
        x"2500",
        x"3230",
        x"2058",
        x"2020",
        x"2020",
        x"0020",
        x"2523",
        x"3230",
        x"2058",
        x"2020",
        x"2020",
        x"2500",
        x"3430",
        x"2058",
        x"2020",
        x"0020",
        x"2041",
        x"2020",
        x"2020",
        x"2020",
        x"2000",
        x"2020",
        x"2020",
        x"2020",
        x"0020",
        x"0020",
        x"6325",
        x"2500",
        x"3430",
        x"2058",
        x"203A",
        x"0000",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"010E",
        x"0C00",
        x"0D0D",
        x"0C00",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0606",
        x"0000",
        x"010E",
        x"0D00",
        x"0D0D",
        x"0000",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0000",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0F00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0606",
        x"0000",
        x"000E",
        x"1000",
        x"0D0D",
        x"0300",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0706",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0400",
        x"0408",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0706",
        x"0000",
        x"000E",
        x"0D00",
        x"0E0D",
        x"0400",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0400",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0B00",
        x"4223",
        x"3C42",
        x"0223",
        x"2542",
        x"0223",
        x"3C42",
        x"0223",
        x"0942",
        x"2323",
        x"3B42",
        x"0223",
        x"0E42",
        x"1923",
        x"3B42",
        x"0223",
        x"1D42",
        x"4201",
        x"0642",
        x"2C01",
        x"2942",
        x"2C01",
        x"0642",
        x"2C01",
        x"0742",
        x"0101",
        x"0642",
        x"2C01",
        x"3142",
        x"1501",
        x"0642",
        x"2C01",
        x"2E42",
        x"4218",
        x"4242",
        x"2118",
        x"2442",
        x"2118",
        x"1C42",
        x"2118",
        x"0C42",
        x"1818",
        x"4242",
        x"2118",
        x"1042",
        x"2718",
        x"4242",
        x"2118",
        x"2F42",
        x"4200",
        x"3842",
        x"2D00",
        x"2842",
        x"2D00",
        x"1C42",
        x"2D00",
        x"0D42",
        x"0000",
        x"3842",
        x"2D00",
        x"3342",
        x"2B00",
        x"1C42",
        x"2D00",
        x"0A42",
        x"4234",
        x"3742",
        x"3634",
        x"1742",
        x"3E06",
        x"3742",
        x"3634",
        x"0342",
        x"3434",
        x"3742",
        x"3634",
        x"4042",
        x"3F34",
        x"3842",
        x"3834",
        x"2042",
        x"1F1E",
        x"2042",
        x"1F1E",
        x"3A42",
        x"391E",
        x"2042",
        x"1F1E",
        x"0442",
        x"1E1E",
        x"2042",
        x"1F1E",
        x"1142",
        x"3D1E",
        x"2042",
        x"1F1E",
        x"1442",
        x"4212",
        x"1442",
        x"1512",
        x"1B42",
        x"1612",
        x"1441",
        x"1512",
        x"0842",
        x"1212",
        x"4242",
        x"1512",
        x"0F42",
        x"2612",
        x"4235",
        x"1512",
        x"1342",
        x"4230",
        x"1342",
        x"1930",
        x"1A42",
        x"2230",
        x"1342",
        x"1930",
        x"0542",
        x"3030",
        x"4242",
        x"1930",
        x"3242",
        x"2A30",
        x"4242",
        x"1930",
        x"4142",
        x"4344",
        x"4E41",
        x"4144",
        x"4C53",
        x"4342",
        x"4243",
        x"5343",
        x"4542",
        x"4251",
        x"5449",
        x"4D42",
        x"4249",
        x"454E",
        x"5042",
        x"424C",
        x"4152",
        x"5242",
        x"424B",
        x"4356",
        x"5642",
        x"4353",
        x"434C",
        x"4C43",
        x"4344",
        x"494C",
        x"4C43",
        x"4356",
        x"504D",
        x"5043",
        x"4358",
        x"5950",
        x"4544",
        x"4443",
        x"5845",
        x"4544",
        x"4559",
        x"524F",
        x"4E49",
        x"4943",
        x"584E",
        x"4E49",
        x"4A59",
        x"504D",
        x"534A",
        x"4C52",
        x"4144",
        x"444C",
        x"4C58",
        x"5944",
        x"534C",
        x"4E52",
        x"504F",
        x"524F",
        x"5041",
        x"4148",
        x"4850",
        x"5050",
        x"5848",
        x"4850",
        x"5059",
        x"414C",
        x"4C50",
        x"5050",
        x"584C",
        x"4C50",
        x"5259",
        x"4C4F",
        x"4F52",
        x"5252",
        x"4954",
        x"5452",
        x"5353",
        x"4342",
        x"4553",
        x"5343",
        x"4445",
        x"4553",
        x"5349",
        x"4154",
        x"5453",
        x"5350",
        x"5854",
        x"5453",
        x"5359",
        x"5A54",
        x"4154",
        x"5458",
        x"5941",
        x"5254",
        x"5442",
        x"4253",
        x"5354",
        x"5458",
        x"4158",
        x"5854",
        x"5453",
        x"4159",
        x"4157",
        x"2D49",
        x"2D2D",
        x"0A00",
        x"2500",
        x"0063",
        x"2020",
        x"7453",
        x"7461",
        x"7375",
        x"203A",
        x"3600",
        x"3035",
        x"2032",
        x"6552",
        x"6967",
        x"7473",
        x"7265",
        x"3A73",
        x"200A",
        x"4120",
        x"253D",
        x"3230",
        x"2058",
        x"3D58",
        x"3025",
        x"5832",
        x"5920",
        x"253D",
        x"3230",
        x"2058",
        x"5053",
        x"303D",
        x"2531",
        x"3230",
        x"2058",
        x"4350",
        x"253D",
        x"3430",
        x"0A58",
        x"0000",
        x"2411",
        x"BE1F",
        x"EFCF",
        x"E0DF",
        x"BFDE",
        x"BFCD",
        x"E013",
        x"E6A0",
        x"E0B0",
        x"E0EA",
        x"E3FC",
        x"EF0F",
        x"9503",
        x"BF0B",
        x"C004",
        x"95D8",
        x"920D",
        x"9631",
        x"F3C8",
        x"34AE",
        x"07B1",
        x"F7C9",
        x"E023",
        x"E4AE",
        x"E0B3",
        x"C001",
        x"921D",
        x"3BA2",
        x"07B2",
        x"F7E1",
        x"940E",
        x"1617",
        x"940C",
        x"1E03",
        x"940C",
        x"0000",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"E68F",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E0C0",
        x"E0D0",
        x"940E",
        x"1409",
        x"2EF8",
        x"E088",
        x"16F8",
        x"F461",
        x"9720",
        x"F3C1",
        x"9721",
        x"940E",
        x"13E8",
        x"E280",
        x"940E",
        x"13E8",
        x"E088",
        x"940E",
        x"13E8",
        x"CFEE",
        x"E08D",
        x"16F8",
        x"F4C1",
        x"9720",
        x"F441",
        x"2FC0",
        x"2FD1",
        x"9189",
        x"2388",
        x"F031",
        x"940E",
        x"13E8",
        x"CFFA",
        x"0FC0",
        x"1FD1",
        x"8218",
        x"E08A",
        x"940E",
        x"13E8",
        x"E08D",
        x"940E",
        x"13E8",
        x"B7CD",
        x"B7DE",
        x"E0E5",
        x"940C",
        x"1692",
        x"E18F",
        x"158F",
        x"F684",
        x"2D8F",
        x"940E",
        x"13E8",
        x"2FE0",
        x"2FF1",
        x"0FEC",
        x"1FFD",
        x"82F0",
        x"9621",
        x"CFC6",
        x"B330",
        x"B328",
        x"7E20",
        x"BB28",
        x"B328",
        x"2B86",
        x"2B97",
        x"2F68",
        x"6260",
        x"2762",
        x"BB68",
        x"B380",
        x"2783",
        x"FF86",
        x"CFFC",
        x"9508",
        x"E060",
        x"E070",
        x"E182",
        x"E090",
        x"940E",
        x"04A1",
        x"9508",
        x"B392",
        x"7C90",
        x"BB92",
        x"B392",
        x"2B89",
        x"BB82",
        x"E085",
        x"958A",
        x"F7F1",
        x"0000",
        x"B181",
        x"E090",
        x"9508",
        x"E060",
        x"E070",
        x"E180",
        x"E090",
        x"940E",
        x"04A1",
        x"E082",
        x"E090",
        x"940E",
        x"04B8",
        x"9508",
        x"E060",
        x"E070",
        x"E181",
        x"E090",
        x"940E",
        x"04A1",
        x"E082",
        x"E090",
        x"940E",
        x"04B8",
        x"9508",
        x"B392",
        x"7C90",
        x"BB92",
        x"B392",
        x"2B89",
        x"BB82",
        x"E085",
        x"958A",
        x"F7F1",
        x"0000",
        x"B181",
        x"9A90",
        x"E095",
        x"959A",
        x"F7F1",
        x"0000",
        x"B121",
        x"E090",
        x"2B92",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2FC6",
        x"2FD7",
        x"161C",
        x"061D",
        x"F464",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E084",
        x"E090",
        x"940E",
        x"04A1",
        x"9516",
        x"9507",
        x"9721",
        x"CFF1",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"2EE6",
        x"2EF7",
        x"2F04",
        x"2F15",
        x"2FC2",
        x"E160",
        x"E070",
        x"940E",
        x"04EF",
        x"E160",
        x"E070",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"04EF",
        x"E06A",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"04EF",
        x"E064",
        x"E070",
        x"2F8C",
        x"E090",
        x"940E",
        x"04EF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"9508",
        x"2F28",
        x"2F39",
        x"5220",
        x"0931",
        x"352F",
        x"0531",
        x"F010",
        x"E28E",
        x"E090",
        x"939F",
        x"938F",
        x"E68C",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FD6",
        x"2FC7",
        x"937F",
        x"936F",
        x"939F",
        x"938F",
        x"E58D",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"2F8D",
        x"2F9C",
        x"940E",
        x"0531",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"E0C8",
        x"E0D0",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E08C",
        x"E090",
        x"940E",
        x"04A1",
        x"9516",
        x"9507",
        x"9721",
        x"F7A1",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"E1C0",
        x"E0D0",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E08C",
        x"E090",
        x"940E",
        x"04A1",
        x"9516",
        x"9507",
        x"9721",
        x"F7A1",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"93CF",
        x"93DF",
        x"E520",
        x"E033",
        x"933F",
        x"932F",
        x"E324",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"0587",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E0CA",
        x"E0D0",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"1428",
        x"9390",
        x"0351",
        x"9380",
        x"0350",
        x"9721",
        x"F7A1",
        x"91DF",
        x"91CF",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"5F2E",
        x"4F3F",
        x"933F",
        x"932F",
        x"E321",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"818B",
        x"819C",
        x"940E",
        x"0587",
        x"808B",
        x"809C",
        x"2CA1",
        x"2CB1",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"8189",
        x"819A",
        x"E0A0",
        x"E0B0",
        x"1588",
        x"0599",
        x"05AA",
        x"05BB",
        x"F11C",
        x"940E",
        x"04D0",
        x"E028",
        x"E030",
        x"0CCC",
        x"1CDD",
        x"1CEE",
        x"1CFF",
        x"2F48",
        x"2F59",
        x"7041",
        x"2755",
        x"E060",
        x"E070",
        x"2AC4",
        x"2AD5",
        x"2AE6",
        x"2AF7",
        x"9596",
        x"9587",
        x"FEE0",
        x"C004",
        x"E24D",
        x"26C4",
        x"24EE",
        x"24FF",
        x"5021",
        x"0931",
        x"F739",
        x"EF8F",
        x"1A88",
        x"0A98",
        x"0AA8",
        x"0AB8",
        x"CFD4",
        x"92FF",
        x"92EF",
        x"92DF",
        x"92CF",
        x"EB80",
        x"E091",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"E060",
        x"E070",
        x"E183",
        x"E090",
        x"940E",
        x"04A1",
        x"9508",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"5F2E",
        x"4F3F",
        x"933F",
        x"932F",
        x"5F2E",
        x"4F3F",
        x"933F",
        x"932F",
        x"E22E",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"818A",
        x"938F",
        x"8189",
        x"938F",
        x"818C",
        x"938F",
        x"818B",
        x"938F",
        x"818E",
        x"938F",
        x"818D",
        x"938F",
        x"EB8B",
        x"E091",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"8189",
        x"819A",
        x"940E",
        x"056E",
        x"818D",
        x"819E",
        x"940E",
        x"0587",
        x"80CD",
        x"80DE",
        x"2CE1",
        x"2CF1",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"818B",
        x"819C",
        x"E0A0",
        x"E0B0",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F044",
        x"940E",
        x"064A",
        x"EF9F",
        x"1AC9",
        x"0AD9",
        x"0AE9",
        x"0AF9",
        x"CFEF",
        x"9626",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"9508",
        x"E060",
        x"E070",
        x"E184",
        x"E090",
        x"940E",
        x"04A1",
        x"E082",
        x"E090",
        x"940E",
        x"04B8",
        x"9508",
        x"E060",
        x"E070",
        x"E185",
        x"E090",
        x"940E",
        x"04A1",
        x"E082",
        x"E090",
        x"940E",
        x"04B8",
        x"9508",
        x"E060",
        x"E070",
        x"E186",
        x"E090",
        x"940E",
        x"04A1",
        x"9508",
        x"E060",
        x"E070",
        x"E187",
        x"E090",
        x"940E",
        x"04A1",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"0587",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1428",
        x"91DF",
        x"91CF",
        x"9508",
        x"E2A2",
        x"E0B0",
        x"EEEE",
        x"E0F6",
        x"940C",
        x"1669",
        x"A37A",
        x"A369",
        x"E520",
        x"E033",
        x"933F",
        x"932F",
        x"E324",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"0587",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2CA1",
        x"2CB1",
        x"2E8C",
        x"2E9D",
        x"E221",
        x"0E82",
        x"1C91",
        x"E104",
        x"E011",
        x"2E20",
        x"2E31",
        x"E48F",
        x"2E48",
        x"E084",
        x"2E58",
        x"E49D",
        x"2E69",
        x"E094",
        x"2E79",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2EE8",
        x"2EF9",
        x"2EC8",
        x"2ED9",
        x"A1E9",
        x"A1FA",
        x"9509",
        x"2DEC",
        x"2DFD",
        x"9381",
        x"9391",
        x"2ECE",
        x"2EDF",
        x"15E8",
        x"05F9",
        x"F7A1",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"0D8A",
        x"1D9B",
        x"939F",
        x"938F",
        x"E587",
        x"E094",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2CCE",
        x"2CDF",
        x"2DEC",
        x"2DFD",
        x"8180",
        x"8191",
        x"E0F2",
        x"0ECF",
        x"1CD1",
        x"939F",
        x"938F",
        x"E581",
        x"E094",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"14C8",
        x"04D9",
        x"F731",
        x"925F",
        x"924F",
        x"923F",
        x"922F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2DEE",
        x"2DFF",
        x"9181",
        x"9191",
        x"2EEE",
        x"2EFF",
        x"940E",
        x"0531",
        x"14E8",
        x"04F9",
        x"F7A9",
        x"927F",
        x"926F",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"E1F0",
        x"0EAF",
        x"1CB1",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"14A1",
        x"E021",
        x"06B2",
        x"F009",
        x"CF94",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"9593",
        x"9390",
        x"0351",
        x"9380",
        x"0350",
        x"96A2",
        x"E1E2",
        x"940C",
        x"1685",
        x"ED60",
        x"E074",
        x"940E",
        x"06E8",
        x"9508",
        x"E0A6",
        x"E0B0",
        x"E9EF",
        x"E0F7",
        x"940C",
        x"1675",
        x"2EE6",
        x"2EF7",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"5F2C",
        x"4F3F",
        x"933F",
        x"932F",
        x"E520",
        x"E033",
        x"933F",
        x"932F",
        x"E327",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"E488",
        x"E094",
        x"939F",
        x"938F",
        x"E104",
        x"E011",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"816D",
        x"817E",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"054D",
        x"E486",
        x"E094",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"818D",
        x"819E",
        x"940E",
        x"056E",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"0587",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"5041",
        x"0951",
        x"0961",
        x"0971",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"1618",
        x"0619",
        x"061A",
        x"061B",
        x"F424",
        x"2DEE",
        x"2DFF",
        x"9509",
        x"CFE7",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"9601",
        x"9390",
        x"0351",
        x"9380",
        x"0350",
        x"9626",
        x"E0E6",
        x"940C",
        x"1691",
        x"EB61",
        x"E074",
        x"940E",
        x"0799",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"E1E9",
        x"E0F8",
        x"940C",
        x"166F",
        x"2EC6",
        x"2ED7",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E520",
        x"E033",
        x"933F",
        x"932F",
        x"E32A",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"0587",
        x"2DEC",
        x"2DFD",
        x"9509",
        x"2F08",
        x"2F19",
        x"E481",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"2EE8",
        x"E081",
        x"2EF8",
        x"92FF",
        x"92EF",
        x"940E",
        x"1718",
        x"2F60",
        x"2F71",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"054D",
        x"E38F",
        x"E094",
        x"939F",
        x"938F",
        x"92FF",
        x"92EF",
        x"940E",
        x"1718",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"E290",
        x"2EA9",
        x"E094",
        x"2EB9",
        x"2C8E",
        x"2C9F",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"5041",
        x"0951",
        x"0961",
        x"0971",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"9702",
        x"05A1",
        x"05B1",
        x"F0D4",
        x"2DEC",
        x"2DFD",
        x"9509",
        x"2EE8",
        x"2EF9",
        x"1708",
        x"0719",
        x"F079",
        x"931F",
        x"930F",
        x"92FF",
        x"938F",
        x"92BF",
        x"92AF",
        x"929F",
        x"928F",
        x"940E",
        x"1718",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2D0E",
        x"2D1F",
        x"CFD2",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"9601",
        x"9390",
        x"0351",
        x"9380",
        x"0350",
        x"9624",
        x"E0EC",
        x"940C",
        x"168B",
        x"EC65",
        x"E074",
        x"940E",
        x"0813",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2F86",
        x"2F97",
        x"940E",
        x"04B8",
        x"2FC8",
        x"2FD9",
        x"2F80",
        x"2F91",
        x"940E",
        x"04DB",
        x"2F48",
        x"2F59",
        x"2F8C",
        x"2F9D",
        x"E0A0",
        x"E0B0",
        x"2FA8",
        x"2FB9",
        x"2799",
        x"2788",
        x"E060",
        x"E070",
        x"2F08",
        x"2F19",
        x"2F2A",
        x"2F3B",
        x"2B04",
        x"2B15",
        x"2B26",
        x"2B37",
        x"2F93",
        x"2F82",
        x"2F71",
        x"2F60",
        x"E420",
        x"E432",
        x"E04F",
        x"E050",
        x"940E",
        x"1637",
        x"939F",
        x"938F",
        x"937F",
        x"936F",
        x"935F",
        x"934F",
        x"933F",
        x"932F",
        x"E182",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"B72D",
        x"B73E",
        x"5F24",
        x"4F3F",
        x"B60F",
        x"94F8",
        x"BF3E",
        x"BE0F",
        x"BF2D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"EFEB",
        x"E0F8",
        x"940C",
        x"166F",
        x"2F08",
        x"2F19",
        x"E83C",
        x"2E83",
        x"E030",
        x"2E93",
        x"EA42",
        x"2EA4",
        x"E040",
        x"2EB4",
        x"E081",
        x"E090",
        x"E05C",
        x"2EE5",
        x"E054",
        x"2EF5",
        x"E1C4",
        x"E0D1",
        x"E06F",
        x"2EC6",
        x"E064",
        x"2ED6",
        x"FF00",
        x"C020",
        x"2B89",
        x"F451",
        x"92DF",
        x"92CF",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2DE8",
        x"2DF9",
        x"8181",
        x"938F",
        x"8180",
        x"938F",
        x"92FF",
        x"92EF",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E080",
        x"E090",
        x"9516",
        x"9507",
        x"E0E2",
        x"0E8E",
        x"1C91",
        x"14A8",
        x"04B9",
        x"F6B1",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"168B",
        x"3180",
        x"F4D8",
        x"2FE8",
        x"E0F0",
        x"0FEE",
        x"1FFF",
        x"59E4",
        x"4FFF",
        x"8181",
        x"938F",
        x"8180",
        x"938F",
        x"E080",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"EE8F",
        x"E093",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E7E2",
        x"E0F9",
        x"940C",
        x"166B",
        x"9180",
        x"0352",
        x"9190",
        x"0353",
        x"2B89",
        x"F409",
        x"C065",
        x"E800",
        x"E013",
        x"E982",
        x"2E88",
        x"E083",
        x"2E98",
        x"EA92",
        x"2EC9",
        x"E093",
        x"2ED9",
        x"E724",
        x"2EE2",
        x"E023",
        x"2EF2",
        x"E03F",
        x"2E43",
        x"E031",
        x"2E53",
        x"E1C4",
        x"E0D1",
        x"E04C",
        x"2E64",
        x"E041",
        x"2E74",
        x"E059",
        x"2EA5",
        x"E051",
        x"2EB5",
        x"2D8E",
        x"2D9F",
        x"5784",
        x"4093",
        x"9120",
        x"0352",
        x"9130",
        x"0353",
        x"1782",
        x"0793",
        x"F00C",
        x"C04B",
        x"2FE0",
        x"2FF1",
        x"8140",
        x"8151",
        x"5F0E",
        x"4F1F",
        x"2DE8",
        x"2DF9",
        x"8120",
        x"8131",
        x"E0F2",
        x"0E8F",
        x"1C91",
        x"935F",
        x"934F",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"925F",
        x"924F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"2DEC",
        x"2DFD",
        x"9181",
        x"9191",
        x"2ECE",
        x"2EDF",
        x"940E",
        x"08F5",
        x"927F",
        x"926F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"2DEE",
        x"2DFF",
        x"9181",
        x"2EEE",
        x"2EFF",
        x"940E",
        x"0940",
        x"92BF",
        x"92AF",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"B78D",
        x"B79E",
        x"9642",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"CFB7",
        x"EF85",
        x"E090",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E1E0",
        x"940C",
        x"1687",
        x"E0A0",
        x"E0B0",
        x"EFE7",
        x"E0F9",
        x"940C",
        x"166F",
        x"E086",
        x"E090",
        x"940E",
        x"04DB",
        x"2EE8",
        x"2EF9",
        x"E088",
        x"E090",
        x"940E",
        x"04DB",
        x"2EA8",
        x"2EB9",
        x"E08A",
        x"E090",
        x"940E",
        x"04B8",
        x"2E88",
        x"2E99",
        x"E08B",
        x"E090",
        x"940E",
        x"04B8",
        x"2EC8",
        x"2ED9",
        x"E021",
        x"22C2",
        x"24DD",
        x"E0C1",
        x"E0D0",
        x"C002",
        x"0FCC",
        x"1FDD",
        x"958A",
        x"F7E2",
        x"2F8C",
        x"2F9D",
        x"7A8A",
        x"7092",
        x"2B89",
        x"F031",
        x"E06E",
        x"E070",
        x"E08C",
        x"E090",
        x"940E",
        x"08A7",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"08F5",
        x"92FF",
        x"92EF",
        x"EE82",
        x"E093",
        x"939F",
        x"938F",
        x"E104",
        x"E011",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"23CC",
        x"F0D9",
        x"2F8C",
        x"2F9D",
        x"7C8C",
        x"2799",
        x"2B89",
        x"F019",
        x"ED89",
        x"E093",
        x"C002",
        x"ED80",
        x"E093",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2D68",
        x"2D79",
        x"2D8A",
        x"2D9B",
        x"940E",
        x"054D",
        x"EC8E",
        x"E093",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"75C5",
        x"27DD",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2BCD",
        x"F051",
        x"E06E",
        x"E070",
        x"E08C",
        x"E090",
        x"940E",
        x"08A7",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"06DB",
        x"2D8C",
        x"2D9D",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"168B",
        x"E080",
        x"E090",
        x"940E",
        x"04DB",
        x"9390",
        x"0351",
        x"9380",
        x"0350",
        x"E063",
        x"E070",
        x"E084",
        x"E090",
        x"940E",
        x"08A7",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"06DB",
        x"9390",
        x"034F",
        x"9380",
        x"034E",
        x"9508",
        x"93CF",
        x"93DF",
        x"E481",
        x"E091",
        x"939F",
        x"938F",
        x"E486",
        x"E091",
        x"939F",
        x"938F",
        x"EA8B",
        x"E093",
        x"939F",
        x"938F",
        x"E1C4",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"E580",
        x"E091",
        x"939F",
        x"938F",
        x"E58C",
        x"E091",
        x"939F",
        x"938F",
        x"E985",
        x"E093",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"921F",
        x"E088",
        x"938F",
        x"E781",
        x"E093",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"B78D",
        x"B79E",
        x"9646",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"940E",
        x"0A94",
        x"E483",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"EDC4",
        x"E0D0",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E30B",
        x"E012",
        x"E184",
        x"2EE8",
        x"E081",
        x"2EF8",
        x"E081",
        x"30C6",
        x"07D8",
        x"F091",
        x"8188",
        x"8199",
        x"9622",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"92FF",
        x"92EF",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"CFEA",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"1691",
        x"9140",
        x"0352",
        x"9150",
        x"0353",
        x"E9E2",
        x"E0F3",
        x"E020",
        x"E030",
        x"1724",
        x"0735",
        x"F444",
        x"9161",
        x"9171",
        x"1768",
        x"0779",
        x"F039",
        x"5F2F",
        x"4F3F",
        x"CFF5",
        x"1784",
        x"0795",
        x"F424",
        x"9508",
        x"2F82",
        x"2F93",
        x"9508",
        x"EF8F",
        x"EF9F",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"E2EA",
        x"E0FB",
        x"940C",
        x"1675",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E324",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"80F9",
        x"80EA",
        x"2D8F",
        x"2D9E",
        x"940E",
        x"0B07",
        x"2F08",
        x"2F19",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"FF97",
        x"C012",
        x"92EF",
        x"92FF",
        x"E48F",
        x"E093",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2F80",
        x"2F91",
        x"9622",
        x"E0E6",
        x"940C",
        x"1691",
        x"E061",
        x"E070",
        x"2B89",
        x"F411",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"04A1",
        x"9508",
        x"9360",
        x"037C",
        x"9370",
        x"037D",
        x"9380",
        x"037E",
        x"9390",
        x"037F",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F0B9",
        x"939F",
        x"938F",
        x"937F",
        x"936F",
        x"E189",
        x"E093",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"9508",
        x"E087",
        x"E093",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"EAE8",
        x"E0FB",
        x"940C",
        x"1679",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E32D",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"8169",
        x"817A",
        x"818B",
        x"819C",
        x"940E",
        x"0B6F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9624",
        x"E0E2",
        x"940C",
        x"1695",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F86",
        x"2F97",
        x"940E",
        x"08F5",
        x"93DF",
        x"93CF",
        x"EF89",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"9508",
        x"9180",
        x"0353",
        x"938F",
        x"9180",
        x"0352",
        x"938F",
        x"ED85",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E0E0",
        x"E0FC",
        x"940C",
        x"1671",
        x"E060",
        x"E070",
        x"E082",
        x"E090",
        x"940E",
        x"04A1",
        x"EA82",
        x"2EE8",
        x"E083",
        x"2EF8",
        x"E890",
        x"2EC9",
        x"E093",
        x"2ED9",
        x"E922",
        x"2EA2",
        x"E023",
        x"2EB2",
        x"E704",
        x"E013",
        x"91C0",
        x"0352",
        x"91D0",
        x"0353",
        x"2F80",
        x"2F91",
        x"5784",
        x"4093",
        x"178C",
        x"079D",
        x"F4D4",
        x"2FE0",
        x"2FF1",
        x"9121",
        x"2F0E",
        x"2F1F",
        x"2DEE",
        x"2DFF",
        x"9141",
        x"9151",
        x"2EEE",
        x"2EFF",
        x"2DEC",
        x"2DFD",
        x"9161",
        x"9171",
        x"2ECE",
        x"2EDF",
        x"2DEA",
        x"2DFB",
        x"9181",
        x"9191",
        x"2EAE",
        x"2EBF",
        x"940E",
        x"050B",
        x"CFDB",
        x"30C8",
        x"05D1",
        x"F45C",
        x"E020",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"050B",
        x"9621",
        x"CFF2",
        x"E061",
        x"E070",
        x"E082",
        x"E090",
        x"940E",
        x"04A1",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"168D",
        x"E0A1",
        x"E0B0",
        x"E5E8",
        x"E0FC",
        x"940C",
        x"1675",
        x"2F08",
        x"2F19",
        x"E18F",
        x"8389",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"939F",
        x"938F",
        x"E685",
        x"E091",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1737",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"8189",
        x"3180",
        x"F198",
        x"ED81",
        x"E090",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"8219",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"EC04",
        x"E010",
        x"E124",
        x"2EE2",
        x"E021",
        x"2EF2",
        x"8189",
        x"3180",
        x"F548",
        x"2FE8",
        x"E0F0",
        x"0FEE",
        x"1FFF",
        x"59E4",
        x"4FFF",
        x"8191",
        x"939F",
        x"8190",
        x"939F",
        x"921F",
        x"938F",
        x"931F",
        x"930F",
        x"92FF",
        x"92EF",
        x"940E",
        x"1718",
        x"8189",
        x"5F8F",
        x"8389",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"CFE2",
        x"2F80",
        x"2F91",
        x"940E",
        x"0B24",
        x"FD97",
        x"C008",
        x"2FE8",
        x"2FF9",
        x"58EC",
        x"4FFC",
        x"8129",
        x"8320",
        x"940E",
        x"0BFA",
        x"9621",
        x"E0E6",
        x"940C",
        x"1691",
        x"930F",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"2FAE",
        x"2FBF",
        x"56AE",
        x"4FBC",
        x"2364",
        x"2375",
        x"936D",
        x"937C",
        x"2FAE",
        x"2FBF",
        x"58A0",
        x"4FBC",
        x"934D",
        x"935C",
        x"55EE",
        x"4FFC",
        x"8331",
        x"8320",
        x"2FE8",
        x"2FF9",
        x"58EC",
        x"4FFC",
        x"8300",
        x"940E",
        x"0BFA",
        x"910F",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"9120",
        x"0352",
        x"9130",
        x"0353",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"2FAE",
        x"2FBF",
        x"56AE",
        x"4FBC",
        x"2FCE",
        x"2FDF",
        x"58C0",
        x"4FDC",
        x"2F0E",
        x"2F1F",
        x"550E",
        x"4F1C",
        x"2F48",
        x"2F59",
        x"584C",
        x"4F5C",
        x"1782",
        x"0793",
        x"F4D4",
        x"9601",
        x"9612",
        x"916D",
        x"917C",
        x"9713",
        x"936D",
        x"937D",
        x"816A",
        x"817B",
        x"9369",
        x"9379",
        x"2FE0",
        x"2FF1",
        x"8162",
        x"8173",
        x"9361",
        x"9371",
        x"2F0E",
        x"2F1F",
        x"2FE4",
        x"2FF5",
        x"8161",
        x"9361",
        x"2F4E",
        x"2F5F",
        x"CFE3",
        x"5021",
        x"0931",
        x"9330",
        x"0353",
        x"9320",
        x"0352",
        x"940E",
        x"0BFA",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"940E",
        x"0B24",
        x"2EE8",
        x"2EF9",
        x"FD97",
        x"C030",
        x"EE8B",
        x"E090",
        x"939F",
        x"938F",
        x"E104",
        x"E011",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"2DCE",
        x"2DDF",
        x"0FCC",
        x"1FDD",
        x"2FEC",
        x"2FFD",
        x"55EE",
        x"4FFC",
        x"8180",
        x"8191",
        x"940E",
        x"08F5",
        x"56CE",
        x"4FDC",
        x"8189",
        x"938F",
        x"8188",
        x"938F",
        x"EE81",
        x"E090",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"0CD7",
        x"B78D",
        x"B79E",
        x"960A",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"1691",
        x"E0A5",
        x"E0B0",
        x"E6E4",
        x"E0FD",
        x"940C",
        x"166D",
        x"2EE6",
        x"2EF7",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"E12F",
        x"832D",
        x"2F2C",
        x"2F3D",
        x"5F2B",
        x"4F3F",
        x"933F",
        x"932F",
        x"5024",
        x"0931",
        x"933F",
        x"932F",
        x"5F2E",
        x"4F3F",
        x"933F",
        x"932F",
        x"E62E",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"9180",
        x"0352",
        x"9190",
        x"0353",
        x"80AB",
        x"80BC",
        x"E9E2",
        x"E0F3",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"E000",
        x"E010",
        x"1708",
        x"0719",
        x"F5DC",
        x"9121",
        x"9131",
        x"152A",
        x"053B",
        x"F599",
        x"2FE0",
        x"2FF1",
        x"0FEE",
        x"1FFF",
        x"55EE",
        x"4FFC",
        x"8180",
        x"8191",
        x"2D2E",
        x"2D3F",
        x"2328",
        x"2339",
        x"2B23",
        x"F0C9",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"08F5",
        x"818C",
        x"938F",
        x"818B",
        x"938F",
        x"EB8F",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C099",
        x"812D",
        x"312F",
        x"F431",
        x"2FE0",
        x"2FF1",
        x"58EC",
        x"4FFC",
        x"8120",
        x"832D",
        x"2AE8",
        x"2AF9",
        x"C063",
        x"5F0F",
        x"4F1F",
        x"CFC2",
        x"1708",
        x"0719",
        x"F009",
        x"C05C",
        x"3008",
        x"0511",
        x"F419",
        x"940E",
        x"0BE3",
        x"C080",
        x"818D",
        x"318F",
        x"F411",
        x"E08F",
        x"838D",
        x"2FE0",
        x"2FF1",
        x"0FEE",
        x"1FFF",
        x"2F6E",
        x"2F7F",
        x"566E",
        x"4F7C",
        x"2F2E",
        x"2F3F",
        x"5820",
        x"4F3C",
        x"2F8E",
        x"2F9F",
        x"558E",
        x"4F9C",
        x"2E68",
        x"2E79",
        x"2FA0",
        x"2FB1",
        x"58AC",
        x"4FBC",
        x"2F80",
        x"2F91",
        x"1618",
        x"0619",
        x"F04C",
        x"5F0F",
        x"4F1F",
        x"9310",
        x"0353",
        x"9300",
        x"0352",
        x"2F08",
        x"2F19",
        x"C02D",
        x"2E88",
        x"2E99",
        x"E0F1",
        x"1A8F",
        x"0891",
        x"2FE6",
        x"2FF7",
        x"90D2",
        x"90C2",
        x"2F4E",
        x"2F5F",
        x"5022",
        x"0931",
        x"E0F2",
        x"1A6F",
        x"0871",
        x"9711",
        x"14AC",
        x"04BD",
        x"F718",
        x"2FE6",
        x"2FF7",
        x"82D1",
        x"82C0",
        x"2FE2",
        x"2FF3",
        x"8180",
        x"8191",
        x"8393",
        x"8382",
        x"2DE6",
        x"2DF7",
        x"8180",
        x"8191",
        x"8393",
        x"8382",
        x"918C",
        x"9611",
        x"938C",
        x"9711",
        x"2F64",
        x"2F75",
        x"2D88",
        x"2D99",
        x"CFC7",
        x"2D6E",
        x"2D7F",
        x"818B",
        x"819C",
        x"940E",
        x"0BC6",
        x"816D",
        x"8149",
        x"815A",
        x"2F80",
        x"2F91",
        x"0F88",
        x"1F99",
        x"2FE8",
        x"2FF9",
        x"56EE",
        x"4FFC",
        x"812B",
        x"813C",
        x"2324",
        x"2335",
        x"8331",
        x"8320",
        x"2FE8",
        x"2FF9",
        x"58E0",
        x"4FFC",
        x"8351",
        x"8340",
        x"2FE8",
        x"2FF9",
        x"55EE",
        x"4FFC",
        x"82F1",
        x"82E0",
        x"2FE0",
        x"2FF1",
        x"58EC",
        x"4FFC",
        x"8360",
        x"940E",
        x"0BFA",
        x"9625",
        x"E0EE",
        x"940C",
        x"1689",
        x"E060",
        x"E071",
        x"940E",
        x"0D5E",
        x"9508",
        x"E060",
        x"E072",
        x"940E",
        x"0D5E",
        x"9508",
        x"E061",
        x"E070",
        x"940E",
        x"0D5E",
        x"9508",
        x"E062",
        x"E070",
        x"940E",
        x"0D5E",
        x"9508",
        x"E064",
        x"E070",
        x"940E",
        x"0D5E",
        x"9508",
        x"E068",
        x"E070",
        x"940E",
        x"0D5E",
        x"9508",
        x"3F6F",
        x"EF2F",
        x"0772",
        x"F419",
        x"FF80",
        x"C028",
        x"C02A",
        x"3F6E",
        x"EF3F",
        x"0773",
        x"F419",
        x"FF80",
        x"C024",
        x"C020",
        x"3F6D",
        x"EF2F",
        x"0772",
        x"F429",
        x"2F69",
        x"2777",
        x"EC33",
        x"2783",
        x"C008",
        x"3F6C",
        x"EF3F",
        x"0773",
        x"F451",
        x"2F69",
        x"2777",
        x"E32C",
        x"2782",
        x"2F26",
        x"2F37",
        x"2728",
        x"2F82",
        x"2F93",
        x"9508",
        x"FF77",
        x"C003",
        x"940E",
        x"16F8",
        x"C002",
        x"2F86",
        x"2F97",
        x"2799",
        x"9508",
        x"EA8A",
        x"E090",
        x"9508",
        x"E585",
        x"E090",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"EBE5",
        x"E0FE",
        x"940C",
        x"1669",
        x"2E28",
        x"2E39",
        x"2F06",
        x"2F17",
        x"2FC4",
        x"2FD5",
        x"2F84",
        x"2F95",
        x"940E",
        x"16FD",
        x"2CC2",
        x"2CD3",
        x"2CE1",
        x"2CF1",
        x"2C8C",
        x"2C9D",
        x"2CAE",
        x"2CBF",
        x"2E40",
        x"2E51",
        x"2C61",
        x"2C71",
        x"1448",
        x"0459",
        x"046A",
        x"047B",
        x"F0A4",
        x"2F6C",
        x"2F7D",
        x"2D88",
        x"2D99",
        x"940E",
        x"0E7B",
        x"940E",
        x"056E",
        x"2D88",
        x"2D99",
        x"940E",
        x"0587",
        x"940E",
        x"064A",
        x"EF8F",
        x"1A88",
        x"0A98",
        x"0AA8",
        x"0AB8",
        x"CFE7",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"16FD",
        x"2D82",
        x"2D93",
        x"940E",
        x"0587",
        x"2C81",
        x"2C91",
        x"E902",
        x"E012",
        x"E134",
        x"2EA3",
        x"E031",
        x"2EB3",
        x"144C",
        x"045D",
        x"046E",
        x"047F",
        x"F164",
        x"940E",
        x"04D0",
        x"2E28",
        x"2E39",
        x"2F6C",
        x"2F7D",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"0E7B",
        x"1628",
        x"0639",
        x"F0C9",
        x"923F",
        x"922F",
        x"939F",
        x"938F",
        x"92FF",
        x"92EF",
        x"92DF",
        x"92CF",
        x"931F",
        x"930F",
        x"92BF",
        x"92AF",
        x"940E",
        x"1718",
        x"EF9F",
        x"1A89",
        x"0A99",
        x"B78D",
        x"B79E",
        x"960C",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"EF9F",
        x"1AC9",
        x"0AD9",
        x"0AE9",
        x"0AF9",
        x"CFCF",
        x"2788",
        x"2799",
        x"1B8C",
        x"0B9D",
        x"FD97",
        x"C006",
        x"3086",
        x"0591",
        x"F02C",
        x"E085",
        x"E090",
        x"C002",
        x"E080",
        x"E090",
        x"0F88",
        x"1F99",
        x"2FE8",
        x"2FF9",
        x"5AE0",
        x"4FFF",
        x"8181",
        x"938F",
        x"8180",
        x"938F",
        x"E882",
        x"E092",
        x"939F",
        x"938F",
        x"E104",
        x"E011",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"FDD7",
        x"C010",
        x"93DF",
        x"93CF",
        x"E78C",
        x"E092",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"1481",
        x"0491",
        x"F099",
        x"929F",
        x"928F",
        x"E687",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C00E",
        x"E58D",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E1E2",
        x"940C",
        x"1685",
        x"E0A6",
        x"E0B0",
        x"E8EE",
        x"E0FF",
        x"940C",
        x"1677",
        x"E92C",
        x"EF3F",
        x"833A",
        x"8329",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"5F2E",
        x"4F3F",
        x"933F",
        x"932F",
        x"5F2E",
        x"4F3F",
        x"933F",
        x"932F",
        x"E729",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"8149",
        x"815A",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"816B",
        x"817C",
        x"818D",
        x"819E",
        x"394C",
        x"EF2F",
        x"0752",
        x"F529",
        x"E545",
        x"E050",
        x"940E",
        x"0EAF",
        x"816B",
        x"817C",
        x"EA4A",
        x"E050",
        x"818D",
        x"819E",
        x"940E",
        x"0EAF",
        x"816B",
        x"817C",
        x"EF4F",
        x"E050",
        x"818D",
        x"819E",
        x"940E",
        x"0EAF",
        x"E000",
        x"E010",
        x"816B",
        x"817C",
        x"2F40",
        x"2F51",
        x"818D",
        x"819E",
        x"940E",
        x"0EAF",
        x"5001",
        x"0911",
        x"3F08",
        x"EF8F",
        x"0718",
        x"F791",
        x"C002",
        x"940E",
        x"0EAF",
        x"9626",
        x"E0E4",
        x"940C",
        x"1693",
        x"93CF",
        x"93DF",
        x"9B87",
        x"C00B",
        x"940E",
        x"09F1",
        x"2FC8",
        x"2FD9",
        x"E060",
        x"E070",
        x"E089",
        x"E090",
        x"940E",
        x"04A1",
        x"C002",
        x"E0C1",
        x"E0D0",
        x"940E",
        x"140F",
        x"2388",
        x"F031",
        x"940E",
        x"1409",
        x"308D",
        x"F411",
        x"E0C0",
        x"E0D0",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"9508",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E32D",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"1618",
        x"0619",
        x"061A",
        x"061B",
        x"F07C",
        x"E183",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C078",
        x"93BF",
        x"93AF",
        x"939F",
        x"938F",
        x"EF88",
        x"E091",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"9040",
        x"037C",
        x"9050",
        x"037D",
        x"9060",
        x"037E",
        x"9070",
        x"037F",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"24CC",
        x"94C3",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"ED04",
        x"E011",
        x"E194",
        x"2EA9",
        x"E091",
        x"2EB9",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F40C",
        x"C048",
        x"E060",
        x"E070",
        x"E088",
        x"E090",
        x"940E",
        x"04A1",
        x"940E",
        x"0FE2",
        x"2B89",
        x"F499",
        x"92FF",
        x"92EF",
        x"92DF",
        x"92CF",
        x"931F",
        x"930F",
        x"92BF",
        x"92AF",
        x"940E",
        x"1718",
        x"80C9",
        x"80DA",
        x"80EB",
        x"80FC",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"16C8",
        x"06D9",
        x"06EA",
        x"06FB",
        x"F091",
        x"9180",
        x"037C",
        x"9190",
        x"037D",
        x"91A0",
        x"037E",
        x"91B0",
        x"037F",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F081",
        x"E091",
        x"1A49",
        x"0851",
        x"0861",
        x"0871",
        x"F451",
        x"940E",
        x"0A7B",
        x"9040",
        x"037C",
        x"9050",
        x"037D",
        x"9060",
        x"037E",
        x"9070",
        x"037F",
        x"EF8F",
        x"1AC8",
        x"0AD8",
        x"0AE8",
        x"0AF8",
        x"CFAE",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"9508",
        x"E48E",
        x"E092",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"E061",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"04A1",
        x"E78B",
        x"E09F",
        x"9701",
        x"F7F1",
        x"C000",
        x"0000",
        x"E060",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"04A1",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"940E",
        x"10D3",
        x"940E",
        x"0A7B",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"EFEF",
        x"E1F0",
        x"940C",
        x"1679",
        x"821A",
        x"8219",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E72F",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"E080",
        x"E090",
        x"940E",
        x"0B64",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"8189",
        x"819A",
        x"2B89",
        x"F011",
        x"940E",
        x"10D3",
        x"EA8F",
        x"E090",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"940E",
        x"0FE2",
        x"2B89",
        x"F7E1",
        x"EA82",
        x"E090",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"E081",
        x"E090",
        x"940E",
        x"0B64",
        x"940E",
        x"0A7B",
        x"9180",
        x"0350",
        x"9190",
        x"0351",
        x"940E",
        x"0B07",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"FD97",
        x"C00C",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"55EE",
        x"4FFC",
        x"8120",
        x"8131",
        x"FF32",
        x"C002",
        x"940E",
        x"0CD7",
        x"9622",
        x"E0E2",
        x"940C",
        x"1695",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"9180",
        x"0352",
        x"9190",
        x"0353",
        x"3088",
        x"0591",
        x"F419",
        x"940E",
        x"0BE3",
        x"C032",
        x"2F28",
        x"2F39",
        x"5F2F",
        x"4F3F",
        x"9330",
        x"0353",
        x"9320",
        x"0352",
        x"2F28",
        x"2F39",
        x"0F22",
        x"1F33",
        x"2FE2",
        x"2FF3",
        x"56EE",
        x"4FFC",
        x"9140",
        x"034E",
        x"9150",
        x"034F",
        x"8351",
        x"8340",
        x"2FE2",
        x"2FF3",
        x"58E0",
        x"4FFC",
        x"EF4F",
        x"EF5F",
        x"8351",
        x"8340",
        x"2FE2",
        x"2FF3",
        x"55EE",
        x"4FFC",
        x"E040",
        x"E055",
        x"8351",
        x"8340",
        x"2FE8",
        x"2FF9",
        x"58EC",
        x"4FFC",
        x"E02F",
        x"8320",
        x"940E",
        x"0BFA",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"10F9",
        x"91DF",
        x"91CF",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"EAE6",
        x"E1F1",
        x"940C",
        x"1679",
        x"940E",
        x"1409",
        x"8389",
        x"940E",
        x"1409",
        x"838A",
        x"2F8C",
        x"2F9D",
        x"9603",
        x"939F",
        x"938F",
        x"E882",
        x"E091",
        x"939F",
        x"938F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"818B",
        x"819C",
        x"9120",
        x"0390",
        x"9130",
        x"0391",
        x"0F28",
        x"1F39",
        x"2733",
        x"9330",
        x"0391",
        x"9320",
        x"0390",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9624",
        x"E0E2",
        x"940C",
        x"1695",
        x"E0A0",
        x"E0B0",
        x"EDE9",
        x"E1F1",
        x"940C",
        x"1669",
        x"E98E",
        x"E091",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"940E",
        x"1409",
        x"2F08",
        x"0F88",
        x"0B11",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2CA1",
        x"2CB1",
        x"24CC",
        x"94CA",
        x"2CDC",
        x"2C71",
        x"2C51",
        x"2CE1",
        x"2CF1",
        x"2C81",
        x"2C91",
        x"3503",
        x"0511",
        x"F191",
        x"EFCF",
        x"EFDF",
        x"940E",
        x"140F",
        x"2388",
        x"F009",
        x"C098",
        x"9721",
        x"F7C9",
        x"92FF",
        x"92EF",
        x"929F",
        x"928F",
        x"E784",
        x"E091",
        x"939F",
        x"938F",
        x"E1C4",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"92BF",
        x"92AF",
        x"92DF",
        x"92CF",
        x"925F",
        x"927F",
        x"E48B",
        x"E091",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"B78D",
        x"B79E",
        x"9642",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"B7CD",
        x"B7DE",
        x"E1E2",
        x"940C",
        x"1685",
        x"940E",
        x"1409",
        x"2F08",
        x"2E08",
        x"0C00",
        x"0B11",
        x"3301",
        x"0511",
        x"F099",
        x"931F",
        x"938F",
        x"E38D",
        x"E091",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"CFAF",
        x"E081",
        x"E090",
        x"9390",
        x"0391",
        x"9380",
        x"0390",
        x"940E",
        x"11A0",
        x"2F08",
        x"2F19",
        x"940E",
        x"11A0",
        x"2FC8",
        x"940E",
        x"11A0",
        x"2E3C",
        x"2C21",
        x"0D82",
        x"1D93",
        x"5003",
        x"0911",
        x"2DC7",
        x"2DD5",
        x"2E68",
        x"2E79",
        x"1A6C",
        x"0A7D",
        x"2C46",
        x"2C57",
        x"0E4C",
        x"1E5D",
        x"1610",
        x"0611",
        x"F4C4",
        x"940E",
        x"11A0",
        x"144C",
        x"045D",
        x"F410",
        x"2CC4",
        x"2CD5",
        x"14A4",
        x"04B5",
        x"F410",
        x"2CA4",
        x"2CB5",
        x"940E",
        x"056E",
        x"2D84",
        x"2D95",
        x"940E",
        x"0587",
        x"940E",
        x"064A",
        x"9621",
        x"5001",
        x"0911",
        x"CFE1",
        x"940E",
        x"11A0",
        x"940E",
        x"1409",
        x"2F08",
        x"0F88",
        x"0B11",
        x"9180",
        x"0390",
        x"9190",
        x"0391",
        x"2B89",
        x"F021",
        x"EF9F",
        x"1AE9",
        x"0AF9",
        x"C003",
        x"EF2F",
        x"1A82",
        x"0A92",
        x"2E7C",
        x"2E5D",
        x"CF5E",
        x"940E",
        x"1409",
        x"2F08",
        x"0F88",
        x"0B11",
        x"CF58",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F06",
        x"2F17",
        x"939F",
        x"938F",
        x"E38A",
        x"E091",
        x"939F",
        x"938F",
        x"E1C4",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2B01",
        x"F019",
        x"E28E",
        x"E091",
        x"C002",
        x"E284",
        x"E091",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"EDE3",
        x"E1F2",
        x"940C",
        x"1679",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E324",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1737",
        x"8189",
        x"819A",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"3084",
        x"0591",
        x"F448",
        x"B328",
        x"732F",
        x"E036",
        x"0F88",
        x"1F99",
        x"953A",
        x"F7E1",
        x"2B82",
        x"BB88",
        x"B368",
        x"7860",
        x"E070",
        x"E886",
        x"E091",
        x"940E",
        x"129F",
        x"B368",
        x"7460",
        x"E070",
        x"E88A",
        x"E091",
        x"940E",
        x"129F",
        x"9622",
        x"E0E2",
        x"940C",
        x"1695",
        x"BA1A",
        x"EF8F",
        x"BB87",
        x"E38F",
        x"BB81",
        x"B812",
        x"BA18",
        x"E020",
        x"EE31",
        x"E040",
        x"E050",
        x"E060",
        x"EE71",
        x"E080",
        x"E090",
        x"940E",
        x"1414",
        x"940E",
        x"0A94",
        x"940E",
        x"0BFA",
        x"E060",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"04A1",
        x"E060",
        x"E070",
        x"E08A",
        x"E090",
        x"940E",
        x"04A1",
        x"E081",
        x"E090",
        x"940E",
        x"0B64",
        x"E061",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"0B6F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E3ED",
        x"E1F3",
        x"940C",
        x"1671",
        x"2EB8",
        x"2EA9",
        x"2F48",
        x"2F59",
        x"2EE4",
        x"2EF5",
        x"1AE8",
        x"0AF9",
        x"2F04",
        x"2F15",
        x"5F4F",
        x"4F5F",
        x"2FE0",
        x"2FF1",
        x"8120",
        x"5621",
        x"312A",
        x"F390",
        x"ED94",
        x"2EC9",
        x"E090",
        x"2ED9",
        x"E0C0",
        x"E0D0",
        x"2DEC",
        x"2DFD",
        x"9181",
        x"9191",
        x"2ECE",
        x"2EDF",
        x"2FE8",
        x"2FF9",
        x"9001",
        x"2000",
        x"F7E9",
        x"9731",
        x"2F4E",
        x"2F5F",
        x"1B48",
        x"0B59",
        x"16E4",
        x"06F5",
        x"F414",
        x"2D4E",
        x"2D5F",
        x"2D6B",
        x"2D7A",
        x"940E",
        x"1708",
        x"2B89",
        x"F451",
        x"0FCC",
        x"1FDD",
        x"55CE",
        x"4FDF",
        x"81E8",
        x"81F9",
        x"2F80",
        x"2F91",
        x"9509",
        x"C016",
        x"9621",
        x"31C9",
        x"05D1",
        x"F6B9",
        x"92AF",
        x"92BF",
        x"E88E",
        x"E090",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"168D",
        x"93CF",
        x"93DF",
        x"E886",
        x"E094",
        x"939F",
        x"938F",
        x"E0C6",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"E78F",
        x"E094",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"9508",
        x"93CF",
        x"93DF",
        x"3081",
        x"F419",
        x"940E",
        x"1395",
        x"C01A",
        x"E78A",
        x"E094",
        x"939F",
        x"938F",
        x"E1C4",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"E783",
        x"E094",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"9508",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"E188",
        x"B98A",
        x"EF67",
        x"E17E",
        x"E08F",
        x"E090",
        x"940E",
        x"1637",
        x"5021",
        x"B929",
        x"9508",
        x"9508",
        x"9B5D",
        x"CFFE",
        x"B98C",
        x"9508",
        x"308D",
        x"F011",
        x"308A",
        x"F439",
        x"3061",
        x"F049",
        x"E08D",
        x"940E",
        x"13E8",
        x"E08A",
        x"C002",
        x"3061",
        x"F011",
        x"940E",
        x"13E8",
        x"9508",
        x"E060",
        x"940E",
        x"13EC",
        x"E080",
        x"E090",
        x"9508",
        x"E061",
        x"940E",
        x"13EC",
        x"E080",
        x"E090",
        x"9508",
        x"9508",
        x"9B5F",
        x"CFFE",
        x"B18C",
        x"9508",
        x"E080",
        x"9508",
        x"B18B",
        x"7880",
        x"9508",
        x"E080",
        x"9508",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F429",
        x"E188",
        x"B98A",
        x"E686",
        x"B989",
        x"C002",
        x"940E",
        x"13D8",
        x"E080",
        x"940E",
        x"13B4",
        x"940E",
        x"1395",
        x"9508",
        x"9508",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E2EE",
        x"E1F4",
        x"940C",
        x"166A",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"04D0",
        x"2F08",
        x"2F19",
        x"2FE8",
        x"2FF9",
        x"5BED",
        x"4FFA",
        x"95C8",
        x"2C30",
        x"2CE3",
        x"2CF1",
        x"E083",
        x"16E8",
        x"04F1",
        x"F06C",
        x"940E",
        x"04D0",
        x"2E78",
        x"2E69",
        x"E09C",
        x"16E9",
        x"04F1",
        x"F03C",
        x"940E",
        x"04D0",
        x"2E58",
        x"2E49",
        x"C004",
        x"2C71",
        x"2C61",
        x"2C51",
        x"2C41",
        x"2FE0",
        x"2FF1",
        x"5BED",
        x"4FF9",
        x"95C8",
        x"2D80",
        x"E090",
        x"E063",
        x"E070",
        x"940E",
        x"1626",
        x"2E88",
        x"2E99",
        x"93DF",
        x"93CF",
        x"E38B",
        x"E095",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E000",
        x"E010",
        x"E398",
        x"2EA9",
        x"E095",
        x"2EB9",
        x"E124",
        x"2EC2",
        x"E021",
        x"2ED2",
        x"2DE8",
        x"2DF9",
        x"0FE0",
        x"1FF1",
        x"5BED",
        x"4FF8",
        x"95C8",
        x"2DE0",
        x"921F",
        x"93EF",
        x"92BF",
        x"92AF",
        x"E184",
        x"2EE8",
        x"E081",
        x"2EF8",
        x"92DF",
        x"92CF",
        x"940E",
        x"1718",
        x"5F0F",
        x"4F1F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"3003",
        x"0511",
        x"F709",
        x"E386",
        x"E095",
        x"939F",
        x"938F",
        x"92FF",
        x"92EF",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2D83",
        x"E090",
        x"3181",
        x"0591",
        x"F008",
        x"C0CD",
        x"2FE8",
        x"2FF9",
        x"5DE0",
        x"4FFF",
        x"940C",
        x"165E",
        x"E28D",
        x"E095",
        x"C002",
        x"E284",
        x"E095",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C0B5",
        x"2F8C",
        x"2F9D",
        x"9602",
        x"0D87",
        x"1D91",
        x"FC77",
        x"959A",
        x"939F",
        x"938F",
        x"E18B",
        x"E095",
        x"C004",
        x"926F",
        x"927F",
        x"E180",
        x"E095",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"9621",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C095",
        x"926F",
        x"927F",
        x"E085",
        x"E095",
        x"CFEB",
        x"926F",
        x"927F",
        x"EF8A",
        x"E094",
        x"CFE6",
        x"926F",
        x"927F",
        x"EE8F",
        x"E094",
        x"CFE1",
        x"926F",
        x"927F",
        x"EE84",
        x"E094",
        x"CFDC",
        x"926F",
        x"927F",
        x"ED89",
        x"E094",
        x"CFD7",
        x"926F",
        x"927F",
        x"EC8E",
        x"E094",
        x"CFD2",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"EC81",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C05F",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"EB84",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C047",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"EA87",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C02F",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"E98A",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C017",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"E88D",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"E88B",
        x"E094",
        x"939F",
        x"938F",
        x"E184",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"B7CD",
        x"B7DE",
        x"E1E1",
        x"940C",
        x"1686",
        x"E0A0",
        x"E0B0",
        x"E9E4",
        x"E1F5",
        x"940C",
        x"1671",
        x"E283",
        x"E090",
        x"940E",
        x"04B8",
        x"2F08",
        x"2F19",
        x"E286",
        x"E090",
        x"940E",
        x"04DB",
        x"2EB8",
        x"2EA9",
        x"E284",
        x"E090",
        x"940E",
        x"04B8",
        x"2ED8",
        x"2EC9",
        x"E282",
        x"E090",
        x"940E",
        x"04B8",
        x"2EF8",
        x"2EE9",
        x"E281",
        x"E090",
        x"940E",
        x"04B8",
        x"2FC8",
        x"2FD9",
        x"E280",
        x"E090",
        x"940E",
        x"04B8",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93DF",
        x"93CF",
        x"939F",
        x"938F",
        x"E18D",
        x"E098",
        x"939F",
        x"938F",
        x"E1C4",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"E182",
        x"E098",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1718",
        x"B78D",
        x"B79E",
        x"9642",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"E2C2",
        x"E0D1",
        x"E02F",
        x"2EC2",
        x"E028",
        x"2ED2",
        x"E134",
        x"2EE3",
        x"E031",
        x"2EF3",
        x"FF07",
        x"C005",
        x"8188",
        x"2E08",
        x"0C00",
        x"0B99",
        x"C002",
        x"E28D",
        x"E090",
        x"939F",
        x"938F",
        x"92DF",
        x"92CF",
        x"E184",
        x"2EA8",
        x"E081",
        x"2EB8",
        x"92FF",
        x"92EF",
        x"940E",
        x"1718",
        x"0F00",
        x"1F11",
        x"9621",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E091",
        x"32CA",
        x"07D9",
        x"F6F1",
        x"E08D",
        x"E098",
        x"939F",
        x"938F",
        x"92BF",
        x"92AF",
        x"940E",
        x"1718",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"168D",
        x"940E",
        x"130B",
        x"E080",
        x"E090",
        x"940E",
        x"10F9",
        x"E584",
        x"E093",
        x"940E",
        x"0450",
        x"E584",
        x"E093",
        x"940E",
        x"1337",
        x"CFF7",
        x"2400",
        x"2755",
        x"C004",
        x"0E08",
        x"1F59",
        x"0F88",
        x"1F99",
        x"9700",
        x"F029",
        x"9576",
        x"9567",
        x"F3B8",
        x"0571",
        x"F7B9",
        x"2D80",
        x"2F95",
        x"9508",
        x"E2A1",
        x"2E1A",
        x"1BAA",
        x"1BBB",
        x"2FEA",
        x"2FFB",
        x"C00D",
        x"1FAA",
        x"1FBB",
        x"1FEE",
        x"1FFF",
        x"17A2",
        x"07B3",
        x"07E4",
        x"07F5",
        x"F020",
        x"1BA2",
        x"0BB3",
        x"0BE4",
        x"0BF5",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"941A",
        x"F769",
        x"9560",
        x"9570",
        x"9580",
        x"9590",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"0FEE",
        x"1FFF",
        x"2400",
        x"1C00",
        x"BE0B",
        x"95D8",
        x"920F",
        x"9631",
        x"95D8",
        x"920F",
        x"9508",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"1BCA",
        x"0BDB",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"9409",
        x"882A",
        x"8839",
        x"8848",
        x"845F",
        x"846E",
        x"847D",
        x"848C",
        x"849B",
        x"84AA",
        x"84B9",
        x"84C8",
        x"80DF",
        x"80EE",
        x"80FD",
        x"810C",
        x"811B",
        x"81AA",
        x"81B9",
        x"0FCE",
        x"1DD1",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2FCA",
        x"2FDB",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"8168",
        x"8179",
        x"818A",
        x"819B",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F421",
        x"E264",
        x"ED79",
        x"E58B",
        x"E097",
        x"E12D",
        x"EF33",
        x"E041",
        x"E050",
        x"940E",
        x"1DE4",
        x"2E82",
        x"2E93",
        x"2EA4",
        x"2EB5",
        x"EA27",
        x"E431",
        x"E040",
        x"E050",
        x"940E",
        x"1DC9",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"EE2C",
        x"EF34",
        x"EF4F",
        x"EF5F",
        x"2D9B",
        x"2D8A",
        x"2D79",
        x"2D68",
        x"940E",
        x"1DC9",
        x"2FB9",
        x"2FA8",
        x"2F97",
        x"2F86",
        x"0D8C",
        x"1D9D",
        x"1DAE",
        x"1DBF",
        x"FFB7",
        x"C003",
        x"9701",
        x"09A1",
        x"48B0",
        x"8388",
        x"8399",
        x"83AA",
        x"83BB",
        x"779F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"940E",
        x"16A1",
        x"9508",
        x"E28A",
        x"E091",
        x"940E",
        x"16A1",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"9380",
        x"012A",
        x"9390",
        x"012B",
        x"93A0",
        x"012C",
        x"93B0",
        x"012D",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"5041",
        x"4050",
        x"F030",
        x"918D",
        x"9001",
        x"1980",
        x"F419",
        x"2000",
        x"F7B9",
        x"1B88",
        x"0B99",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E1EE",
        x"E1F7",
        x"940C",
        x"1677",
        x"810F",
        x"8518",
        x"2FE0",
        x"2FF1",
        x"8183",
        x"6088",
        x"8383",
        x"2F4C",
        x"2F5D",
        x"5F45",
        x"4F5F",
        x"8569",
        x"857A",
        x"2F80",
        x"2F91",
        x"940E",
        x"1752",
        x"2FE0",
        x"2FF1",
        x"8123",
        x"7F27",
        x"8323",
        x"E0E4",
        x"940C",
        x"1693",
        x"E0AE",
        x"E0B0",
        x"E3ED",
        x"E1F7",
        x"940C",
        x"1679",
        x"E085",
        x"838C",
        x"898B",
        x"899C",
        x"839A",
        x"8389",
        x"2F4C",
        x"2F5D",
        x"5E49",
        x"4F5F",
        x"896D",
        x"897E",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"1B41",
        x"962E",
        x"E0E2",
        x"940C",
        x"1695",
        x"E0AB",
        x"E0B0",
        x"E5E8",
        x"E1F7",
        x"940C",
        x"1669",
        x"2EC8",
        x"2ED9",
        x"2EE6",
        x"2EF7",
        x"2F04",
        x"2F15",
        x"2FE8",
        x"2FF9",
        x"8217",
        x"8216",
        x"8183",
        x"FF81",
        x"C1FF",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2E68",
        x"2E79",
        x"2DEC",
        x"2DFD",
        x"8193",
        x"2DEE",
        x"2DFF",
        x"FD93",
        x"95C8",
        x"FF93",
        x"8000",
        x"9631",
        x"2D80",
        x"2EEE",
        x"2EFF",
        x"2388",
        x"F409",
        x"C1E5",
        x"3285",
        x"F451",
        x"FD93",
        x"95C8",
        x"FF93",
        x"8000",
        x"9631",
        x"2D80",
        x"2EEE",
        x"2EFF",
        x"3285",
        x"F431",
        x"2D6C",
        x"2D7D",
        x"E090",
        x"940E",
        x"1CFC",
        x"CFDE",
        x"2C91",
        x"2C21",
        x"2C31",
        x"E1FF",
        x"15F3",
        x"F0E0",
        x"328B",
        x"F079",
        x"F438",
        x"3280",
        x"F079",
        x"3283",
        x"F4A9",
        x"2D23",
        x"6120",
        x"C010",
        x"328D",
        x"F059",
        x"3380",
        x"F471",
        x"2D23",
        x"6021",
        x"C009",
        x"2D83",
        x"6082",
        x"2E38",
        x"2DE3",
        x"60E4",
        x"C024",
        x"2DF3",
        x"60F8",
        x"C027",
        x"2E32",
        x"C029",
        x"FC37",
        x"C034",
        x"ED20",
        x"0F28",
        x"302A",
        x"F498",
        x"FE36",
        x"C007",
        x"2D89",
        x"E06A",
        x"940E",
        x"1DC0",
        x"2E92",
        x"0E98",
        x"C01A",
        x"2D82",
        x"E06A",
        x"940E",
        x"1DC0",
        x"2E22",
        x"0E28",
        x"2D83",
        x"6280",
        x"2E38",
        x"C010",
        x"328E",
        x"F431",
        x"FC36",
        x"C194",
        x"2DE3",
        x"64E0",
        x"2E3E",
        x"C008",
        x"368C",
        x"F421",
        x"2DF3",
        x"68F0",
        x"2E3F",
        x"C002",
        x"3688",
        x"F469",
        x"2DEE",
        x"2DFF",
        x"FD93",
        x"95C8",
        x"FF93",
        x"8000",
        x"9631",
        x"2D80",
        x"2EEE",
        x"2EFF",
        x"2388",
        x"F009",
        x"CFAB",
        x"2F98",
        x"7D9F",
        x"5495",
        x"3093",
        x"F428",
        x"5F0C",
        x"4F1F",
        x"E32F",
        x"8329",
        x"C00E",
        x"3683",
        x"F031",
        x"3783",
        x"F081",
        x"3583",
        x"F009",
        x"C06B",
        x"C028",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"8389",
        x"5F0E",
        x"4F1F",
        x"2488",
        x"9483",
        x"2C91",
        x"2CA6",
        x"2CB7",
        x"C018",
        x"2E40",
        x"2E51",
        x"E0F2",
        x"0E4F",
        x"1C51",
        x"2FE0",
        x"2FF1",
        x"80A0",
        x"80B1",
        x"FE36",
        x"C003",
        x"2D69",
        x"E070",
        x"C002",
        x"EF6F",
        x"EF7F",
        x"2D8A",
        x"2D9B",
        x"940E",
        x"1CB1",
        x"2E88",
        x"2E99",
        x"2D04",
        x"2D15",
        x"2DF3",
        x"77FF",
        x"2E3F",
        x"C01B",
        x"2E40",
        x"2E51",
        x"E022",
        x"0E42",
        x"1C51",
        x"2FE0",
        x"2FF1",
        x"80A0",
        x"80B1",
        x"FE36",
        x"C003",
        x"2D69",
        x"E070",
        x"C002",
        x"EF6F",
        x"EF7F",
        x"2D8A",
        x"2D9B",
        x"940E",
        x"1CA4",
        x"2E88",
        x"2E99",
        x"2DF3",
        x"68F0",
        x"2E3F",
        x"2D04",
        x"2D15",
        x"FC33",
        x"C021",
        x"2D82",
        x"E090",
        x"1688",
        x"0699",
        x"F4E0",
        x"2D6C",
        x"2D7D",
        x"E280",
        x"E090",
        x"940E",
        x"1CFC",
        x"942A",
        x"CFF3",
        x"2DEA",
        x"2DFB",
        x"FC37",
        x"95C8",
        x"FE37",
        x"8000",
        x"9631",
        x"2D80",
        x"2EAE",
        x"2EBF",
        x"2D6C",
        x"2D7D",
        x"E090",
        x"940E",
        x"1CFC",
        x"1021",
        x"942A",
        x"E021",
        x"1A82",
        x"0891",
        x"1481",
        x"0491",
        x"F749",
        x"C0F4",
        x"3684",
        x"F011",
        x"3689",
        x"F551",
        x"2FE0",
        x"2FF1",
        x"FE37",
        x"C007",
        x"8160",
        x"8171",
        x"8182",
        x"8193",
        x"5F0C",
        x"4F1F",
        x"C008",
        x"8160",
        x"8171",
        x"2E07",
        x"0C00",
        x"0B88",
        x"0B99",
        x"5F0E",
        x"4F1F",
        x"2DF3",
        x"76FF",
        x"2E3F",
        x"FF97",
        x"C009",
        x"9590",
        x"9580",
        x"9570",
        x"9561",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"68F0",
        x"2E3F",
        x"E02A",
        x"E030",
        x"2D46",
        x"2D57",
        x"940E",
        x"1D59",
        x"2E88",
        x"1886",
        x"C047",
        x"3785",
        x"F431",
        x"2D23",
        x"7E2F",
        x"2EB2",
        x"E02A",
        x"E030",
        x"C025",
        x"2D93",
        x"7F99",
        x"2EB9",
        x"368F",
        x"F0C1",
        x"F418",
        x"3588",
        x"F079",
        x"C0C0",
        x"3780",
        x"F019",
        x"3788",
        x"F021",
        x"C0BB",
        x"2FE9",
        x"61E0",
        x"2EBE",
        x"FEB4",
        x"C00D",
        x"2DFB",
        x"60F4",
        x"2EBF",
        x"C009",
        x"FE34",
        x"C00A",
        x"2F29",
        x"6026",
        x"2EB2",
        x"C006",
        x"E028",
        x"E030",
        x"C005",
        x"E120",
        x"E030",
        x"C002",
        x"E120",
        x"E032",
        x"2FE0",
        x"2FF1",
        x"FEB7",
        x"C007",
        x"8160",
        x"8171",
        x"8182",
        x"8193",
        x"5F0C",
        x"4F1F",
        x"C006",
        x"8160",
        x"8171",
        x"E080",
        x"E090",
        x"5F0E",
        x"4F1F",
        x"2D46",
        x"2D57",
        x"940E",
        x"1D59",
        x"2E88",
        x"1886",
        x"2DFB",
        x"77FF",
        x"2E3F",
        x"FE36",
        x"C00D",
        x"2D23",
        x"7F2E",
        x"2EA2",
        x"1489",
        x"F458",
        x"FE34",
        x"C00B",
        x"FC32",
        x"C009",
        x"2D83",
        x"7E8E",
        x"2EA8",
        x"C005",
        x"2CB8",
        x"2CA3",
        x"C003",
        x"2CB8",
        x"C001",
        x"2CB9",
        x"FEA4",
        x"C010",
        x"2FEC",
        x"2FFD",
        x"0DE8",
        x"1DF1",
        x"8180",
        x"3380",
        x"F421",
        x"2D9A",
        x"7E99",
        x"2EA9",
        x"C009",
        x"FEA2",
        x"C006",
        x"94B3",
        x"94B3",
        x"C004",
        x"2D8A",
        x"7886",
        x"F009",
        x"94B3",
        x"FCA3",
        x"C012",
        x"FEA0",
        x"C006",
        x"14B2",
        x"F490",
        x"0C28",
        x"2C92",
        x"189B",
        x"C00F",
        x"14B2",
        x"F468",
        x"2D6C",
        x"2D7D",
        x"E280",
        x"E090",
        x"940E",
        x"1CFC",
        x"94B3",
        x"CFF6",
        x"14B2",
        x"F418",
        x"182B",
        x"C002",
        x"2C98",
        x"2C21",
        x"FEA4",
        x"C012",
        x"2D6C",
        x"2D7D",
        x"E380",
        x"E090",
        x"940E",
        x"1CFC",
        x"FEA2",
        x"C019",
        x"FCA1",
        x"C003",
        x"E788",
        x"E090",
        x"C002",
        x"E588",
        x"E090",
        x"2D6C",
        x"2D7D",
        x"C00D",
        x"2D8A",
        x"7886",
        x"F061",
        x"FEA1",
        x"C002",
        x"E28B",
        x"C001",
        x"E280",
        x"FCA7",
        x"E28D",
        x"2D6C",
        x"2D7D",
        x"E090",
        x"940E",
        x"1CFC",
        x"1489",
        x"F440",
        x"2D6C",
        x"2D7D",
        x"E380",
        x"E090",
        x"940E",
        x"1CFC",
        x"949A",
        x"CFF6",
        x"948A",
        x"2DE6",
        x"2DF7",
        x"0DE8",
        x"1DF1",
        x"8180",
        x"2D6C",
        x"2D7D",
        x"E090",
        x"940E",
        x"1CFC",
        x"2088",
        x"F799",
        x"2022",
        x"F409",
        x"CE13",
        x"2D6C",
        x"2D7D",
        x"E280",
        x"E090",
        x"940E",
        x"1CFC",
        x"942A",
        x"CFF5",
        x"2DEC",
        x"2DFD",
        x"8186",
        x"8197",
        x"C002",
        x"EF8F",
        x"EF9F",
        x"962B",
        x"E1E2",
        x"940C",
        x"1685",
        x"FD20",
        x"C00A",
        x"2FE8",
        x"2FF9",
        x"FD23",
        x"C005",
        x"FF22",
        x"C002",
        x"8373",
        x"8362",
        x"8351",
        x"8340",
        x"9508",
        x"FD44",
        x"C01D",
        x"FD46",
        x"C01D",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"2FA4",
        x"2FB5",
        x"2FE6",
        x"2FF7",
        x"0FAA",
        x"1FBB",
        x"1FEE",
        x"1FFF",
        x"9410",
        x"F7D1",
        x"0F4A",
        x"1F5B",
        x"1F6E",
        x"1F7F",
        x"2F97",
        x"2F86",
        x"2F75",
        x"2F64",
        x"0F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"C009",
        x"E033",
        x"C001",
        x"E034",
        x"0F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"5031",
        x"F7D1",
        x"0F62",
        x"1D71",
        x"1D81",
        x"1D91",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2F80",
        x"2F91",
        x"940E",
        x"1CBD",
        x"2FC8",
        x"2FD9",
        x"FD97",
        x"C00A",
        x"940E",
        x"1C8C",
        x"2B89",
        x"F7A1",
        x"2F60",
        x"2F71",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1D3F",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2FD6",
        x"2EE4",
        x"2EF5",
        x"2EB2",
        x"940E",
        x"1CBD",
        x"2F28",
        x"2F39",
        x"2733",
        x"322B",
        x"0531",
        x"F031",
        x"322D",
        x"0531",
        x"F469",
        x"2D8B",
        x"6880",
        x"2EB8",
        x"50D1",
        x"F411",
        x"E080",
        x"C077",
        x"2F80",
        x"2F91",
        x"940E",
        x"1CBD",
        x"FD97",
        x"CFF8",
        x"2DCB",
        x"7FCD",
        x"2D2B",
        x"7320",
        x"F521",
        x"3380",
        x"F511",
        x"24AA",
        x"94AA",
        x"0EAD",
        x"F409",
        x"C04D",
        x"2F80",
        x"2F91",
        x"940E",
        x"1CBD",
        x"FD97",
        x"C047",
        x"2F28",
        x"2F39",
        x"7D2F",
        x"2733",
        x"3528",
        x"0531",
        x"F451",
        x"64C2",
        x"50D2",
        x"F1E9",
        x"2F80",
        x"2F91",
        x"940E",
        x"1CBD",
        x"FF97",
        x"C007",
        x"C036",
        x"FEB6",
        x"C002",
        x"60C2",
        x"C001",
        x"61C2",
        x"2DDA",
        x"2C81",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"ED20",
        x"0F28",
        x"3028",
        x"F088",
        x"FFC4",
        x"C005",
        x"2F60",
        x"2F71",
        x"940E",
        x"1D3F",
        x"C01E",
        x"302A",
        x"F040",
        x"FFC6",
        x"CFF7",
        x"7D2F",
        x"EE3F",
        x"0F32",
        x"3036",
        x"F790",
        x"5027",
        x"2F4C",
        x"2D9B",
        x"2D8A",
        x"2D79",
        x"2D68",
        x"940E",
        x"1977",
        x"2E86",
        x"2E97",
        x"2EA8",
        x"2EB9",
        x"60C2",
        x"50D1",
        x"F069",
        x"2F80",
        x"2F91",
        x"940E",
        x"1CBD",
        x"FF97",
        x"CFD7",
        x"FDC1",
        x"C005",
        x"CF9F",
        x"2C81",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"FFC7",
        x"C008",
        x"94B0",
        x"94A0",
        x"9490",
        x"9480",
        x"1C81",
        x"1C91",
        x"1CA1",
        x"1CB1",
        x"2F2C",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"196A",
        x"E081",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"E2A0",
        x"E0B0",
        x"E6ED",
        x"E1FA",
        x"940C",
        x"166C",
        x"2EA8",
        x"2EB9",
        x"2E96",
        x"2EE4",
        x"2EF5",
        x"2FE2",
        x"2FF3",
        x"2F0C",
        x"2F1D",
        x"5F0F",
        x"4F1F",
        x"2EC0",
        x"2ED1",
        x"E280",
        x"2FA0",
        x"2FB1",
        x"921D",
        x"958A",
        x"F7E9",
        x"2DAA",
        x"2DBB",
        x"9613",
        x"908C",
        x"E080",
        x"E090",
        x"2C61",
        x"2C71",
        x"E030",
        x"E061",
        x"E070",
        x"FC83",
        x"95C8",
        x"FE83",
        x"8000",
        x"9631",
        x"2D20",
        x"2F0E",
        x"2F1F",
        x"2E52",
        x"2322",
        x"F419",
        x"E080",
        x"E090",
        x"C0A4",
        x"352E",
        x"F411",
        x"9700",
        x"F169",
        x"2F43",
        x"E050",
        x"1748",
        x"0759",
        x"F43C",
        x"352D",
        x"F171",
        x"322D",
        x"F419",
        x"2077",
        x"F121",
        x"C003",
        x"2077",
        x"F409",
        x"C079",
        x"2D45",
        x"9546",
        x"9546",
        x"9546",
        x"2DAC",
        x"2DBD",
        x"0FA4",
        x"1DB1",
        x"2D45",
        x"7047",
        x"2F06",
        x"2F17",
        x"C002",
        x"0F00",
        x"1F11",
        x"954A",
        x"F7E2",
        x"2F40",
        x"2F51",
        x"915C",
        x"2B45",
        x"934C",
        x"1465",
        x"F059",
        x"1456",
        x"F410",
        x"9453",
        x"CFE4",
        x"945A",
        x"CFE2",
        x"E031",
        x"C004",
        x"2477",
        x"9473",
        x"C001",
        x"2C71",
        x"9601",
        x"CFB9",
        x"2077",
        x"F019",
        x"818E",
        x"6280",
        x"838E",
        x"2333",
        x"F419",
        x"2488",
        x"9483",
        x"C01C",
        x"2DEC",
        x"2DFD",
        x"2F2C",
        x"2F3D",
        x"5D2F",
        x"4F3F",
        x"8180",
        x"9580",
        x"9381",
        x"172E",
        x"073F",
        x"F7D1",
        x"CFF0",
        x"14E1",
        x"04F1",
        x"F041",
        x"2DAE",
        x"2DBF",
        x"938C",
        x"2DEE",
        x"2DFF",
        x"9631",
        x"2EEE",
        x"2EFF",
        x"949A",
        x"2C81",
        x"2099",
        x"F121",
        x"2D8A",
        x"2D9B",
        x"940E",
        x"1CBD",
        x"FD97",
        x"C01B",
        x"2FE8",
        x"2FF9",
        x"27FF",
        x"E023",
        x"95F5",
        x"95E7",
        x"952A",
        x"F7E1",
        x"0DEC",
        x"1DFD",
        x"8120",
        x"E030",
        x"2F48",
        x"2F59",
        x"7047",
        x"2755",
        x"C002",
        x"9535",
        x"9527",
        x"954A",
        x"F7E2",
        x"FD20",
        x"CFD4",
        x"2D6A",
        x"2D7B",
        x"940E",
        x"1D3F",
        x"2088",
        x"F009",
        x"CF7A",
        x"14E1",
        x"04F1",
        x"F019",
        x"2DAE",
        x"2DBF",
        x"921C",
        x"2F80",
        x"2F91",
        x"C018",
        x"2F42",
        x"9546",
        x"9546",
        x"9546",
        x"2DAC",
        x"2DBD",
        x"0FA4",
        x"1DB1",
        x"2F42",
        x"7047",
        x"2F06",
        x"2F17",
        x"C002",
        x"0F00",
        x"1F11",
        x"954A",
        x"F7E2",
        x"2F40",
        x"2F51",
        x"915C",
        x"2B45",
        x"934C",
        x"2E62",
        x"CF93",
        x"96A0",
        x"E0EF",
        x"940C",
        x"1688",
        x"E0A0",
        x"E0B0",
        x"E4E7",
        x"E1FB",
        x"940C",
        x"166C",
        x"2EC8",
        x"2ED9",
        x"2FC6",
        x"2FD7",
        x"2EA4",
        x"2EB5",
        x"2FE8",
        x"2FF9",
        x"8217",
        x"8216",
        x"2C51",
        x"2DEC",
        x"2DFD",
        x"80E3",
        x"2FEC",
        x"2FFD",
        x"FCE3",
        x"95C8",
        x"FEE3",
        x"8000",
        x"9631",
        x"2D80",
        x"2F18",
        x"2FCE",
        x"2FDF",
        x"2388",
        x"F409",
        x"C11F",
        x"E090",
        x"940E",
        x"1C8C",
        x"2B89",
        x"F029",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"19A4",
        x"CFE5",
        x"3215",
        x"F461",
        x"2FEC",
        x"2FFD",
        x"FCE3",
        x"95C8",
        x"FEE3",
        x"8000",
        x"9631",
        x"2D10",
        x"2FCE",
        x"2FDF",
        x"3215",
        x"F4A1",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"1CBD",
        x"FD97",
        x"C0FF",
        x"2F41",
        x"E050",
        x"2F28",
        x"2F39",
        x"2733",
        x"1724",
        x"0735",
        x"F409",
        x"CFC8",
        x"2D6C",
        x"2D7D",
        x"940E",
        x"1D3F",
        x"C0F3",
        x"321A",
        x"F451",
        x"FCE3",
        x"95C8",
        x"FEE3",
        x"8000",
        x"9631",
        x"2D10",
        x"2FCE",
        x"2FDF",
        x"E001",
        x"C001",
        x"E000",
        x"2CF1",
        x"ED20",
        x"0F21",
        x"302A",
        x"F4A0",
        x"6002",
        x"2D6F",
        x"E070",
        x"E080",
        x"E090",
        x"E240",
        x"940E",
        x"1977",
        x"2EF6",
        x"2FEC",
        x"2FFD",
        x"FCE3",
        x"95C8",
        x"FEE3",
        x"8000",
        x"9631",
        x"2D10",
        x"2FCE",
        x"2FDF",
        x"CFE8",
        x"FF01",
        x"C003",
        x"20FF",
        x"F419",
        x"C0C8",
        x"24FF",
        x"94FA",
        x"3618",
        x"F019",
        x"361C",
        x"F071",
        x"C018",
        x"2FEC",
        x"2FFD",
        x"FCE3",
        x"95C8",
        x"FEE3",
        x"8000",
        x"9631",
        x"2D10",
        x"2FCE",
        x"2FDF",
        x"3618",
        x"F461",
        x"6008",
        x"6004",
        x"2FEC",
        x"2FFD",
        x"FCE3",
        x"95C8",
        x"FEE3",
        x"8000",
        x"9631",
        x"2D10",
        x"2FCE",
        x"2FDF",
        x"2311",
        x"F409",
        x"C0A6",
        x"2F61",
        x"E070",
        x"E882",
        x"E090",
        x"940E",
        x"1C95",
        x"2B89",
        x"F409",
        x"C09D",
        x"FD00",
        x"C00A",
        x"2DEA",
        x"2DFB",
        x"8080",
        x"8091",
        x"2D8A",
        x"2D9B",
        x"9602",
        x"2EA8",
        x"2EB9",
        x"C002",
        x"2C81",
        x"2C91",
        x"361E",
        x"F461",
        x"2DEC",
        x"2DFD",
        x"8146",
        x"8157",
        x"E060",
        x"E070",
        x"2F20",
        x"2D88",
        x"2D99",
        x"940E",
        x"196A",
        x"CF51",
        x"3613",
        x"F4C9",
        x"FD01",
        x"C002",
        x"24FF",
        x"94F3",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"1CBD",
        x"FD97",
        x"C073",
        x"1481",
        x"0491",
        x"F041",
        x"2DE8",
        x"2DF9",
        x"8380",
        x"2D88",
        x"2D99",
        x"9601",
        x"2E88",
        x"2E99",
        x"94FA",
        x"20FF",
        x"F761",
        x"C060",
        x"351B",
        x"F479",
        x"2F2C",
        x"2F3D",
        x"2D48",
        x"2D59",
        x"2D6F",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"1A67",
        x"2FC8",
        x"2FD9",
        x"2B89",
        x"F009",
        x"C050",
        x"C049",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"19A4",
        x"FD97",
        x"C04D",
        x"361F",
        x"F1A1",
        x"F428",
        x"3614",
        x"F179",
        x"3619",
        x"F191",
        x"C030",
        x"3713",
        x"F089",
        x"3715",
        x"F141",
        x"C02B",
        x"1481",
        x"0491",
        x"F041",
        x"2DE8",
        x"2DF9",
        x"8260",
        x"2D88",
        x"2D99",
        x"9601",
        x"2E88",
        x"2E99",
        x"94FA",
        x"20FF",
        x"F091",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"1CBD",
        x"2E68",
        x"2E79",
        x"FD97",
        x"C00A",
        x"940E",
        x"1C8C",
        x"2B89",
        x"F331",
        x"2D6C",
        x"2D7D",
        x"2D86",
        x"2D97",
        x"940E",
        x"1D3F",
        x"1481",
        x"0491",
        x"F0C9",
        x"2DE8",
        x"2DF9",
        x"8210",
        x"C015",
        x"6200",
        x"C003",
        x"6100",
        x"C001",
        x"6400",
        x"2F20",
        x"2D48",
        x"2D59",
        x"2D6F",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"19C3",
        x"2388",
        x"F431",
        x"2DEC",
        x"2DFD",
        x"8183",
        x"7380",
        x"F429",
        x"C006",
        x"FD00",
        x"CED4",
        x"9453",
        x"CED2",
        x"2055",
        x"F019",
        x"2D85",
        x"E090",
        x"C002",
        x"EF8F",
        x"EF9F",
        x"B7CD",
        x"B7DE",
        x"E0EF",
        x"940C",
        x"1688",
        x"1191",
        x"940C",
        x"1DBD",
        x"3280",
        x"F019",
        x"5089",
        x"5085",
        x"F7C8",
        x"9508",
        x"2FE8",
        x"2FF9",
        x"95C8",
        x"9631",
        x"1606",
        x"F029",
        x"2000",
        x"F7D1",
        x"2D80",
        x"2D91",
        x"9508",
        x"9731",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"2FE8",
        x"2FF9",
        x"95C8",
        x"9631",
        x"5061",
        x"4070",
        x"1001",
        x"F7D0",
        x"9580",
        x"9590",
        x"0F8E",
        x"1F9F",
        x"9508",
        x"2FE8",
        x"2FF9",
        x"5061",
        x"4070",
        x"9001",
        x"1001",
        x"F7D8",
        x"9580",
        x"9590",
        x"0F8E",
        x"1F9F",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"812B",
        x"FF20",
        x"C033",
        x"FF26",
        x"C00A",
        x"7B2F",
        x"832B",
        x"818E",
        x"819F",
        x"9601",
        x"839F",
        x"838E",
        x"818A",
        x"E090",
        x"C029",
        x"FF22",
        x"C00F",
        x"81E8",
        x"81F9",
        x"8180",
        x"2E08",
        x"0C00",
        x"0B99",
        x"9700",
        x"F419",
        x"6220",
        x"832B",
        x"C01A",
        x"9631",
        x"83F9",
        x"83E8",
        x"C00E",
        x"85EA",
        x"85FB",
        x"9509",
        x"FF97",
        x"C009",
        x"812B",
        x"9601",
        x"F011",
        x"E280",
        x"C001",
        x"E180",
        x"2B82",
        x"838B",
        x"C008",
        x"812E",
        x"813F",
        x"5F2F",
        x"4F3F",
        x"833F",
        x"832E",
        x"2799",
        x"C002",
        x"EF8F",
        x"EF9F",
        x"91DF",
        x"91CF",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FE6",
        x"2FF7",
        x"8123",
        x"FD21",
        x"C003",
        x"EF8F",
        x"EF9F",
        x"C032",
        x"FF22",
        x"C017",
        x"8146",
        x"8157",
        x"8124",
        x"8135",
        x"1742",
        x"0753",
        x"F44C",
        x"81A0",
        x"81B1",
        x"2F2A",
        x"2F3B",
        x"5F2F",
        x"4F3F",
        x"8331",
        x"8320",
        x"938C",
        x"8126",
        x"8137",
        x"5F2F",
        x"4F3F",
        x"8337",
        x"8326",
        x"C019",
        x"2F06",
        x"2F17",
        x"2FD9",
        x"2FC8",
        x"2FE6",
        x"2FF7",
        x"8400",
        x"85F1",
        x"2DE0",
        x"9509",
        x"2B89",
        x"F6C1",
        x"2FA0",
        x"2FB1",
        x"9616",
        x"918D",
        x"919C",
        x"9717",
        x"9601",
        x"9617",
        x"939C",
        x"938E",
        x"9716",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"8123",
        x"FF20",
        x"C012",
        x"FD26",
        x"C010",
        x"3F8F",
        x"EF3F",
        x"0793",
        x"F061",
        x"8382",
        x"7D2F",
        x"6420",
        x"8323",
        x"8126",
        x"8137",
        x"5021",
        x"0931",
        x"8337",
        x"8326",
        x"2799",
        x"9508",
        x"EF8F",
        x"EF9F",
        x"9508",
        x"2FE4",
        x"2FF5",
        x"27AA",
        x"3028",
        x"F169",
        x"3120",
        x"F199",
        x"94E8",
        x"936F",
        x"7F6E",
        x"5F6E",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"4FAF",
        x"E0B1",
        x"D041",
        x"E0B4",
        x"D03F",
        x"0F67",
        x"1F78",
        x"1F89",
        x"1F9A",
        x"1DA1",
        x"0F68",
        x"1F79",
        x"1F8A",
        x"1D91",
        x"1DA1",
        x"0F6A",
        x"1D71",
        x"1D81",
        x"1D91",
        x"1DA1",
        x"D023",
        x"F409",
        x"9468",
        x"913F",
        x"2E06",
        x"0C00",
        x"1930",
        x"0C00",
        x"0C00",
        x"1930",
        x"5D30",
        x"9331",
        x"F6CE",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"2F46",
        x"7047",
        x"5D40",
        x"9341",
        x"E0B3",
        x"D00F",
        x"F7C9",
        x"CFF5",
        x"2F46",
        x"704F",
        x"5D40",
        x"334A",
        x"F018",
        x"5D49",
        x"FD31",
        x"5240",
        x"9341",
        x"D002",
        x"F7A9",
        x"CFE9",
        x"E0B4",
        x"95A6",
        x"9597",
        x"9587",
        x"9577",
        x"9567",
        x"95BA",
        x"F7C9",
        x"9700",
        x"0561",
        x"0571",
        x"9508",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"2E0A",
        x"9406",
        x"9557",
        x"9547",
        x"9537",
        x"9527",
        x"95BA",
        x"F7C9",
        x"0F62",
        x"1F73",
        x"1F84",
        x"1F95",
        x"1DA0",
        x"9508",
        x"2799",
        x"2788",
        x"9508",
        x"2400",
        x"FD80",
        x"0E06",
        x"0F66",
        x"F011",
        x"9586",
        x"F7D1",
        x"2D80",
        x"9508",
        x"27EE",
        x"27FF",
        x"27AA",
        x"27BB",
        x"C008",
        x"0FA2",
        x"1FB3",
        x"1FE4",
        x"1FF5",
        x"0F22",
        x"1F33",
        x"1F44",
        x"1F55",
        x"9596",
        x"9587",
        x"9577",
        x"9567",
        x"F398",
        x"4070",
        x"F7A9",
        x"9700",
        x"F799",
        x"2F6A",
        x"2F7B",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"2E05",
        x"FB97",
        x"F41E",
        x"9400",
        x"940E",
        x"1DFB",
        x"FD57",
        x"D007",
        x"940E",
        x"1637",
        x"FC07",
        x"D003",
        x"F44E",
        x"940C",
        x"1DFB",
        x"9550",
        x"9540",
        x"9530",
        x"9521",
        x"4F3F",
        x"4F4F",
        x"4F5F",
        x"9508",
        x"9590",
        x"9580",
        x"9570",
        x"9561",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"9508",
        x"94F8",
        x"CFFF",
        x"018E",
        x"0194",
        x"01A1",
        x"01B6",
        x"01C6",
        x"01DE",
        x"01E5",
        x"01EB",
        x"01EC",
        x"01F3",
        x"01F7",
        x"0202",
        x"0206",
        x"0210",
        x"01F8",
        x"021B",
        x"0203",
        x"0211",
        x"01FF",
        x"0226",
        x"0227",
        x"0230",
        x"0237",
        x"0244",
        x"0251",
        x"025E",
        x"026B",
        x"0277",
        x"0283",
        x"028F",
        x"029B",
        x"02A4",
        x"02AD",
        x"0ACE",
        x"10F9",
        x"115D",
        x"1002",
        x"158E",
        x"05A0",
        x"0651",
        x"05CB",
        x"0794",
        x"08A2",
        x"080E",
        x"0F88",
        x"11D3",
        x"12CD",
        x"10F4",
        x"0BA2",
        x"096C",
        x"0E5D",
        x"0E62",
        x"0E67",
        x"0E6C",
        x"0E71",
        x"0E76",
        x"0D1D",
        x"0C52",
        x"02B7",
        x"02BC",
        x"02C5",
        x"02CA",
        x"02CF",
        x"02D4",
        x"02D8",
        x"02DD",
        x"02E1",
        x"02E5",
        x"02E9",
        x"02ED",
        x"02F2",
        x"02F7",
        x"02FF",
        x"0305",
        x"030B",
        x"0311",
        x"0318",
        x"031F",
        x"0327",
        x"032F",
        x"0337",
        x"033F",
        x"0345",
        x"0000",
        x"0200",
        x"0000",
        x"0000",
        x"1402",
        x"0000",
        x"0000",
        x"0000",
        x"0200",
        x"0000",
        x"0000",
        x"13FC",
        x"0000",
        x"0000",
        x"564E",
        x"422D",
        x"4944",
        x"435A",
        x"0001",
        x"0000",
        x"7825",
        x"2520",
        x"2078",
        x"7825",
        x"2500",
        x"2078",
        x"7825",
        x"2520",
        x"646C",
        x"3000",
        x"392E",
        x"0030",
        x"4349",
        x"2D45",
        x"3536",
        x"3043",
        x"0032",
        x"6F4E",
        x"2076",
        x"3420",
        x"3220",
        x"3130",
        x"0039",
        x"3531",
        x"343A",
        x"3A36",
        x"3531",
        x"2500",
        x"782A",
        x"2520",
        x"6868",
        x"0078",
        x"7825",
        x"2520",
        x"2078",
        x"6825",
        x"7868",
        x"2500",
        x"2078",
        x"7825",
        x"2520",
        x"0064",
        x"3225",
        x"0078",
        x"4D4E",
        x"0049",
        x"5249",
        x"0051",
        x"6946",
        x"6578",
        x"0064",
        x"6843",
        x"6365",
        x"656B",
        x"6272",
        x"616F",
        x"6472",
        x"4900",
        x"766E",
        x"7265",
        x"6573",
        x"6320",
        x"6568",
        x"6B63",
        x"7265",
        x"6F62",
        x"7261",
        x"0064",
        x"6441",
        x"7264",
        x"7365",
        x"2073",
        x"6170",
        x"7474",
        x"7265",
        x"006E",
        x"6E49",
        x"6576",
        x"7372",
        x"2065",
        x"6461",
        x"7264",
        x"7365",
        x"2073",
        x"6170",
        x"7474",
        x"7265",
        x"006E",
        x"6152",
        x"646E",
        x"6D6F",
        x"4E00",
        x"7665",
        x"7265",
        x"7E00",
        x"3054",
        x"6120",
        x"646E",
        x"7E20",
        x"3154",
        x"7E00",
        x"3054",
        x"6120",
        x"646E",
        x"5420",
        x"0031",
        x"547E",
        x"0030",
        x"3054",
        x"7820",
        x"726F",
        x"5420",
        x"0031",
        x"547E",
        x"2030",
        x"726F",
        x"7E20",
        x"3154",
        x"5400",
        x"2030",
        x"6E78",
        x"726F",
        x"5420",
        x"0031",
        x"547E",
        x"2030",
        x"726F",
        x"5420",
        x"0031",
        x"6C41",
        x"6177",
        x"7379",
        x"4D00",
        x"6D65",
        x"5220",
        x"2064",
        x"7242",
        x"706B",
        x"0074",
        x"654D",
        x"206D",
        x"6452",
        x"5720",
        x"7461",
        x"6863",
        x"4D00",
        x"6D65",
        x"5720",
        x"2072",
        x"7242",
        x"706B",
        x"0074",
        x"654D",
        x"206D",
        x"7257",
        x"5720",
        x"7461",
        x"6863",
        x"4900",
        x"204F",
        x"6452",
        x"4220",
        x"6B72",
        x"7470",
        x"4900",
        x"204F",
        x"6452",
        x"5720",
        x"7461",
        x"6863",
        x"4900",
        x"204F",
        x"7257",
        x"4220",
        x"6B72",
        x"7470",
        x"4900",
        x"204F",
        x"7257",
        x"5720",
        x"7461",
        x"6863",
        x"4500",
        x"2078",
        x"7242",
        x"706B",
        x"0074",
        x"7845",
        x"5720",
        x"7461",
        x"6863",
        x"5400",
        x"6172",
        x"736E",
        x"6569",
        x"746E",
        x"6800",
        x"6C65",
        x"0070",
        x"6F63",
        x"746E",
        x"6E69",
        x"6575",
        x"6E00",
        x"7865",
        x"0074",
        x"7473",
        x"7065",
        x"7200",
        x"6765",
        x"0073",
        x"6964",
        x"0073",
        x"6966",
        x"6C6C",
        x"6300",
        x"6372",
        x"6D00",
        x"6D65",
        x"7200",
        x"6D64",
        x"7700",
        x"6D72",
        x"7400",
        x"7365",
        x"0074",
        x"7273",
        x"6365",
        x"7300",
        x"6570",
        x"6963",
        x"6C61",
        x"7200",
        x"7365",
        x"7465",
        x"7400",
        x"6172",
        x"6563",
        x"6200",
        x"696C",
        x"7473",
        x"6200",
        x"6572",
        x"6B61",
        x"0078",
        x"6177",
        x"6374",
        x"7868",
        x"6200",
        x"6572",
        x"6B61",
        x"6D72",
        x"7700",
        x"7461",
        x"6863",
        x"6D72",
        x"6200",
        x"6572",
        x"6B61",
        x"6D77",
        x"7700",
        x"7461",
        x"6863",
        x"6D77",
        x"6300",
        x"656C",
        x"7261",
        x"7400",
        x"6972",
        x"6767",
        x"7265",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000"
    );

begin

    process (cp2)
    begin
        if rising_edge(cp2) then
            if ce = '1' then
                if (we = '1') then
                    RAM(conv_integer(address)) <= din;
                end if;
                dout <= RAM(conv_integer(address));
            end if;
        end if;
    end process;

end RTL;
