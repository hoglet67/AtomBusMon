library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- This contains 0.72 of the ICE T65 (a.k.a AtomCpuMon) firmware

-- For f_log2 definition
use WORK.SynthCtrlPack.all;

entity XPM is
    generic (
        WIDTH : integer;
        SIZE  : integer
    );
    port(
        cp2     : in  std_logic;
        ce      : in  std_logic;
        address : in  std_logic_vector(f_log2(SIZE) - 1 downto 0);
        din     : in  std_logic_vector(WIDTH - 1 downto 0);
        dout    : out std_logic_vector(WIDTH - 1 downto 0);
        we      : in  std_logic
    );
end;

architecture RTL of XPM is
    
    type ram_type is array (0 to SIZE - 1) of std_logic_vector (WIDTH - 1 downto 0);

    signal RAM : ram_type := (
        x"940C",
        x"03FD",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"940C",
        x"041F",
        x"1287",
        x"128A",
        x"134F",
        x"1299",
        x"12A6",
        x"12BA",
        x"12BF",
        x"12C4",
        x"12CE",
        x"12D3",
        x"12C9",
        x"134F",
        x"12D8",
        x"12F0",
        x"1308",
        x"1320",
        x"1338",
        x"6E55",
        x"6E6B",
        x"776F",
        x"206E",
        x"6F63",
        x"6D6D",
        x"6E61",
        x"2064",
        x"7325",
        x"000A",
        x"6E49",
        x"6574",
        x"7272",
        x"7075",
        x"6574",
        x"0A64",
        x"4300",
        x"5550",
        x"6620",
        x"6572",
        x"2065",
        x"7572",
        x"6E6E",
        x"6E69",
        x"2E67",
        x"2E2E",
        x"000A",
        x"6552",
        x"6573",
        x"7474",
        x"6E69",
        x"2067",
        x"5043",
        x"0A55",
        x"4900",
        x"6C6C",
        x"6765",
        x"6C61",
        x"7420",
        x"6972",
        x"6767",
        x"7265",
        x"6320",
        x"646F",
        x"2065",
        x"7328",
        x"6565",
        x"6820",
        x"6C65",
        x"2070",
        x"6F66",
        x"2072",
        x"7274",
        x"6769",
        x"6567",
        x"2072",
        x"6F63",
        x"6564",
        x"2973",
        x"000A",
        x"2020",
        x"2020",
        x"5825",
        x"3D20",
        x"2520",
        x"0A73",
        x"5400",
        x"6972",
        x"6767",
        x"7265",
        x"4320",
        x"646F",
        x"7365",
        x"0A3A",
        x"2000",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"5200",
        x"6D65",
        x"766F",
        x"6E69",
        x"2067",
        x"4E00",
        x"206F",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"6573",
        x"0A74",
        x"2900",
        x"000A",
        x"2820",
        x"2500",
        x"3A64",
        x"2520",
        x"3430",
        x"2058",
        x"616D",
        x"6B73",
        x"2520",
        x"3430",
        x"3A58",
        x"0020",
        x"7263",
        x"3A63",
        x"2520",
        x"3430",
        x"0A58",
        x"5700",
        x"3A72",
        x"2520",
        x"3430",
        x"2058",
        x"6F74",
        x"2520",
        x"3430",
        x"2058",
        x"203D",
        x"3025",
        x"5832",
        x"000A",
        x"6552",
        x"6573",
        x"7474",
        x"6E69",
        x"2067",
        x"5043",
        x"0A55",
        x"5300",
        x"6574",
        x"7070",
        x"6E69",
        x"2067",
        x"6C25",
        x"2064",
        x"6E69",
        x"7473",
        x"7572",
        x"7463",
        x"6F69",
        x"736E",
        x"000A",
        x"754E",
        x"626D",
        x"7265",
        x"6F20",
        x"2066",
        x"6E69",
        x"7473",
        x"6375",
        x"6974",
        x"6E6F",
        x"2073",
        x"756D",
        x"7473",
        x"6220",
        x"2065",
        x"6F70",
        x"6973",
        x"6974",
        x"6576",
        x"000A",
        x"2020",
        x"2020",
        x"7325",
        x"000A",
        x"6F43",
        x"6D6D",
        x"6E61",
        x"7364",
        x"0A3A",
        x"3A00",
        x"7020",
        x"7361",
        x"6573",
        x"0A64",
        x"3A00",
        x"6620",
        x"6961",
        x"656C",
        x"3A64",
        x"2520",
        x"2064",
        x"7265",
        x"6F72",
        x"7372",
        x"000A",
        x"2520",
        x"3230",
        x"0058",
        x"654D",
        x"6F6D",
        x"7972",
        x"7420",
        x"7365",
        x"3A74",
        x"2520",
        x"0073",
        x"6146",
        x"6C69",
        x"6120",
        x"2074",
        x"3025",
        x"6C34",
        x"2058",
        x"5728",
        x"6F72",
        x"6574",
        x"203A",
        x"3025",
        x"5832",
        x"202C",
        x"6552",
        x"6461",
        x"6220",
        x"6361",
        x"206B",
        x"3025",
        x"5832",
        x"0A29",
        x"4100",
        x"6C6C",
        x"2520",
        x"2064",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"7261",
        x"2065",
        x"6C61",
        x"6572",
        x"6461",
        x"2079",
        x"6573",
        x"0A74",
        x"2000",
        x"6C61",
        x"6572",
        x"6461",
        x"2079",
        x"6573",
        x"2074",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"2000",
        x"6573",
        x"2074",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"5400",
        x"6172",
        x"6963",
        x"676E",
        x"6420",
        x"7369",
        x"6261",
        x"656C",
        x"0A64",
        x"5400",
        x"6172",
        x"6963",
        x"676E",
        x"6520",
        x"6576",
        x"7972",
        x"2520",
        x"646C",
        x"6920",
        x"736E",
        x"7274",
        x"6375",
        x"6974",
        x"6E6F",
        x"2073",
        x"6877",
        x"6C69",
        x"2065",
        x"6973",
        x"676E",
        x"656C",
        x"7320",
        x"6574",
        x"7070",
        x"6E69",
        x"0A67",
        x"4200",
        x"6572",
        x"6B61",
        x"6F70",
        x"6E69",
        x"2F74",
        x"6177",
        x"6374",
        x"2068",
        x"6F6E",
        x"2074",
        x"6573",
        x"2074",
        x"7461",
        x"2520",
        x"3430",
        x"0A58",
        x"2500",
        x"2064",
        x"6177",
        x"6374",
        x"6568",
        x"2F73",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"6D69",
        x"6C70",
        x"6D65",
        x"6E65",
        x"6574",
        x"0A64",
        x"4300",
        x"6D6F",
        x"6970",
        x"656C",
        x"2064",
        x"7461",
        x"2520",
        x"2073",
        x"6E6F",
        x"2520",
        x"0A73",
        x"2500",
        x"2073",
        x"6E49",
        x"432D",
        x"7269",
        x"7563",
        x"7469",
        x"4520",
        x"756D",
        x"616C",
        x"6F74",
        x"2072",
        x"6576",
        x"7372",
        x"6F69",
        x"206E",
        x"7325",
        x"000A",
        x"000A",
        x"2520",
        x"3430",
        x"2058",
        x"203D",
        x"3025",
        x"5832",
        x"000A",
        x"7220",
        x"6165",
        x"6964",
        x"676E",
        x"2000",
        x"7277",
        x"7469",
        x"6E69",
        x"0067",
        x"6820",
        x"7469",
        x"6120",
        x"2074",
        x"3025",
        x"5834",
        x"7400",
        x"6972",
        x"6767",
        x"7265",
        x"203A",
        x"4C49",
        x"454C",
        x"4147",
        x"004C",
        x"7274",
        x"6769",
        x"6567",
        x"3A72",
        x"2520",
        x"0073",
        x"7325",
        x"2C00",
        x"0020",
        x"3025",
        x"6C32",
        x"2E64",
        x"3025",
        x"6C36",
        x"3A64",
        x"0020",
        x"6E49",
        x"6F63",
        x"736E",
        x"7369",
        x"6574",
        x"746E",
        x"5220",
        x"3A64",
        x"2520",
        x"3230",
        x"2058",
        x"3E3C",
        x"2520",
        x"3230",
        x"0A58",
        x"5200",
        x"3A64",
        x"2520",
        x"3430",
        x"2058",
        x"203D",
        x"3025",
        x"5832",
        x"000A",
        x"7257",
        x"203A",
        x"3025",
        x"5834",
        x"3D20",
        x"2520",
        x"3230",
        x"0A58",
        x"0A00",
        x"2500",
        x"0063",
        x"0020",
        x"3025",
        x"5832",
        x"0020",
        x"3025",
        x"5834",
        x"0020",
        x"3E3E",
        x"0020",
        x"000A",
        x"2528",
        x"3230",
        x"2558",
        x"3230",
        x"2C58",
        x"2958",
        x"2800",
        x"3025",
        x"5832",
        x"3025",
        x"5832",
        x"2029",
        x"0020",
        x"3025",
        x"5832",
        x"3025",
        x"5832",
        x"592C",
        x"2020",
        x"2500",
        x"3230",
        x"2558",
        x"3230",
        x"2C58",
        x"2058",
        x"0020",
        x"3025",
        x"5832",
        x"3025",
        x"5832",
        x"2020",
        x"2020",
        x"2800",
        x"3025",
        x"5832",
        x"2C29",
        x"2059",
        x"0020",
        x"2528",
        x"3230",
        x"2C58",
        x"2958",
        x"2020",
        x"2800",
        x"3025",
        x"5832",
        x"2029",
        x"2020",
        x"0020",
        x"3025",
        x"5832",
        x"592C",
        x"2020",
        x"2020",
        x"2500",
        x"3230",
        x"2C58",
        x"2058",
        x"2020",
        x"0020",
        x"3025",
        x"5832",
        x"2020",
        x"2020",
        x"2020",
        x"2300",
        x"3025",
        x"5832",
        x"2020",
        x"2020",
        x"0020",
        x"3025",
        x"5834",
        x"2020",
        x"2020",
        x"4100",
        x"2020",
        x"2020",
        x"2020",
        x"0020",
        x"2020",
        x"2020",
        x"2020",
        x"2020",
        x"2000",
        x"2500",
        x"0063",
        x"3025",
        x"5834",
        x"3A20",
        x"0020",
        x"0800",
        x"0000",
        x"0505",
        x"0005",
        x"0400",
        x"0001",
        x"0C0C",
        x"000C",
        x"0903",
        x"000A",
        x"0605",
        x"0006",
        x"0E00",
        x"0001",
        x"0D0C",
        x"000D",
        x"080C",
        x"0000",
        x"0505",
        x"0005",
        x"0400",
        x"0001",
        x"0C0C",
        x"000C",
        x"0903",
        x"000A",
        x"0606",
        x"0006",
        x"0E00",
        x"0001",
        x"0D0D",
        x"000D",
        x"0800",
        x"0000",
        x"0505",
        x"0005",
        x"0400",
        x"0001",
        x"0C0C",
        x"000C",
        x"0903",
        x"000A",
        x"0605",
        x"0006",
        x"0E00",
        x"0000",
        x"0D0C",
        x"000D",
        x"0800",
        x"0000",
        x"0505",
        x"0005",
        x"0400",
        x"0001",
        x"0C0F",
        x"000C",
        x"0903",
        x"000A",
        x"0606",
        x"0006",
        x"0E00",
        x"0000",
        x"0D10",
        x"000D",
        x"0803",
        x"0000",
        x"0505",
        x"0005",
        x"0400",
        x"0000",
        x"0C0C",
        x"000C",
        x"0903",
        x"000A",
        x"0606",
        x"0007",
        x"0E00",
        x"0000",
        x"0D0C",
        x"000D",
        x"0804",
        x"0004",
        x"0505",
        x"0005",
        x"0400",
        x"0000",
        x"0C0C",
        x"000C",
        x"0903",
        x"000A",
        x"0606",
        x"0007",
        x"0E00",
        x"0000",
        x"0D0D",
        x"000E",
        x"0804",
        x"0000",
        x"0505",
        x"0005",
        x"0400",
        x"0000",
        x"0C0C",
        x"000C",
        x"0903",
        x"000A",
        x"0605",
        x"0006",
        x"0E00",
        x"0000",
        x"0D0C",
        x"000D",
        x"0804",
        x"0000",
        x"0505",
        x"0005",
        x"0400",
        x"0000",
        x"0C0C",
        x"000C",
        x"0903",
        x"000A",
        x"0605",
        x"0006",
        x"0E00",
        x"0000",
        x"0D0C",
        x"000D",
        x"230B",
        x"4242",
        x"233C",
        x"4202",
        x"2325",
        x"4202",
        x"233C",
        x"4202",
        x"2309",
        x"4223",
        x"233B",
        x"4202",
        x"230E",
        x"4219",
        x"233B",
        x"4202",
        x"011D",
        x"4242",
        x"0106",
        x"422C",
        x"0129",
        x"422C",
        x"0106",
        x"422C",
        x"0107",
        x"4201",
        x"0106",
        x"422C",
        x"0131",
        x"4215",
        x"0106",
        x"422C",
        x"182E",
        x"4242",
        x"1842",
        x"4221",
        x"1824",
        x"4221",
        x"181C",
        x"4221",
        x"180C",
        x"4218",
        x"1842",
        x"4221",
        x"1810",
        x"4227",
        x"1842",
        x"4221",
        x"002F",
        x"4242",
        x"0038",
        x"422D",
        x"0028",
        x"422D",
        x"001C",
        x"422D",
        x"000D",
        x"4200",
        x"0038",
        x"422D",
        x"0033",
        x"422B",
        x"001C",
        x"422D",
        x"340A",
        x"4242",
        x"3437",
        x"4236",
        x"0617",
        x"423E",
        x"3437",
        x"4236",
        x"3403",
        x"4234",
        x"3437",
        x"4236",
        x"3440",
        x"423F",
        x"3438",
        x"4238",
        x"1E20",
        x"421F",
        x"1E20",
        x"421F",
        x"1E3A",
        x"4239",
        x"1E20",
        x"421F",
        x"1E04",
        x"421E",
        x"1E20",
        x"421F",
        x"1E11",
        x"423D",
        x"1E20",
        x"421F",
        x"1214",
        x"4242",
        x"1214",
        x"4215",
        x"121B",
        x"4116",
        x"1214",
        x"4215",
        x"1208",
        x"4212",
        x"1242",
        x"4215",
        x"120F",
        x"3526",
        x"1242",
        x"4215",
        x"3013",
        x"4242",
        x"3013",
        x"4219",
        x"301A",
        x"4222",
        x"3013",
        x"4219",
        x"3005",
        x"4230",
        x"3042",
        x"4219",
        x"3032",
        x"422A",
        x"3042",
        x"4219",
        x"4441",
        x"4143",
        x"444E",
        x"5341",
        x"424C",
        x"4343",
        x"4342",
        x"4253",
        x"5145",
        x"4942",
        x"4254",
        x"494D",
        x"4E42",
        x"4245",
        x"4C50",
        x"5242",
        x"4241",
        x"4B52",
        x"5642",
        x"4243",
        x"5356",
        x"4C43",
        x"4343",
        x"444C",
        x"4C43",
        x"4349",
        x"564C",
        x"4D43",
        x"4350",
        x"5850",
        x"5043",
        x"4459",
        x"4345",
        x"4544",
        x"4458",
        x"5945",
        x"4F45",
        x"4952",
        x"434E",
        x"4E49",
        x"4958",
        x"594E",
        x"4D4A",
        x"4A50",
        x"5253",
        x"444C",
        x"4C41",
        x"5844",
        x"444C",
        x"4C59",
        x"5253",
        x"4F4E",
        x"4F50",
        x"4152",
        x"4850",
        x"5041",
        x"5048",
        x"4850",
        x"5058",
        x"5948",
        x"4C50",
        x"5041",
        x"504C",
        x"4C50",
        x"5058",
        x"594C",
        x"4F52",
        x"524C",
        x"524F",
        x"5452",
        x"5249",
        x"5354",
        x"4253",
        x"5343",
        x"4345",
        x"4553",
        x"5344",
        x"4945",
        x"5453",
        x"5341",
        x"5054",
        x"5453",
        x"5358",
        x"5954",
        x"5453",
        x"545A",
        x"5841",
        x"4154",
        x"5459",
        x"4252",
        x"5354",
        x"5442",
        x"5853",
        x"5854",
        x"5441",
        x"5358",
        x"5954",
        x"5741",
        x"4941",
        x"2D2D",
        x"002D",
        x"000A",
        x"6325",
        x"2000",
        x"5320",
        x"6174",
        x"7574",
        x"3A73",
        x"0020",
        x"3536",
        x"3230",
        x"5220",
        x"6765",
        x"7369",
        x"6574",
        x"7372",
        x"0A3A",
        x"2020",
        x"3D41",
        x"3025",
        x"5832",
        x"5820",
        x"253D",
        x"3230",
        x"2058",
        x"3D59",
        x"3025",
        x"5832",
        x"5320",
        x"3D50",
        x"3025",
        x"5834",
        x"5020",
        x"3D43",
        x"3025",
        x"5834",
        x"000A",
        x"5B1B",
        x"3B30",
        x"4830",
        x"1B00",
        x"325B",
        x"004A",
        x"5B1B",
        x"3B30",
        x"4830",
        x"1B00",
        x"325B",
        x"004A",
        x"6463",
        x"6E69",
        x"706F",
        x"7573",
        x"5878",
        x"005B",
        x"2411",
        x"BE1F",
        x"EFCF",
        x"E0DF",
        x"BFDE",
        x"BFCD",
        x"E013",
        x"E6A0",
        x"E0B0",
        x"E0EE",
        x"E3F9",
        x"EF0F",
        x"9503",
        x"BF0B",
        x"C004",
        x"95D8",
        x"920D",
        x"9631",
        x"F3C8",
        x"30AC",
        x"07B1",
        x"F7C9",
        x"E013",
        x"E0AC",
        x"E0B3",
        x"C001",
        x"921D",
        x"37A4",
        x"07B1",
        x"F7E1",
        x"940E",
        x"1481",
        x"940C",
        x"1C85",
        x"940C",
        x"0000",
        x"E0A1",
        x"E0B0",
        x"E2E7",
        x"E0F4",
        x"940C",
        x"14D4",
        x"2F08",
        x"2F19",
        x"E088",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2CE1",
        x"2CF1",
        x"940E",
        x"1462",
        x"2F98",
        x"3088",
        x"F481",
        x"14E1",
        x"04F1",
        x"F3C1",
        x"E081",
        x"1AE8",
        x"08F1",
        x"E088",
        x"940E",
        x"1441",
        x"E280",
        x"940E",
        x"1441",
        x"E088",
        x"940E",
        x"1441",
        x"CFEB",
        x"308D",
        x"F4E1",
        x"14E1",
        x"04F1",
        x"F451",
        x"2FA0",
        x"2FB1",
        x"918D",
        x"2F0A",
        x"2F1B",
        x"2388",
        x"F041",
        x"940E",
        x"1441",
        x"CFF6",
        x"2DEE",
        x"2DFF",
        x"0FE0",
        x"1FF1",
        x"8210",
        x"E08A",
        x"940E",
        x"1441",
        x"E08D",
        x"940E",
        x"1441",
        x"9621",
        x"E0E6",
        x"940C",
        x"14F0",
        x"3280",
        x"F25C",
        x"8399",
        x"940E",
        x"1441",
        x"2FE0",
        x"2FF1",
        x"0DEE",
        x"1DFF",
        x"8199",
        x"8390",
        x"EFBF",
        x"1AEB",
        x"0AFB",
        x"CFBE",
        x"B328",
        x"7C20",
        x"BB28",
        x"B328",
        x"2B68",
        x"2B79",
        x"2B26",
        x"BB28",
        x"E08A",
        x"958A",
        x"F7F1",
        x"C000",
        x"9AC5",
        x"E08A",
        x"958A",
        x"F7F1",
        x"C000",
        x"9508",
        x"E060",
        x"E070",
        x"E182",
        x"E090",
        x"940E",
        x"047B",
        x"9508",
        x"B392",
        x"7C90",
        x"BB92",
        x"B392",
        x"2B98",
        x"BB92",
        x"E085",
        x"958A",
        x"F7F1",
        x"0000",
        x"B181",
        x"E090",
        x"9508",
        x"E060",
        x"E070",
        x"E180",
        x"E090",
        x"940E",
        x"047B",
        x"E385",
        x"958A",
        x"F7F1",
        x"E082",
        x"E090",
        x"940E",
        x"0494",
        x"9508",
        x"E060",
        x"E070",
        x"E181",
        x"E090",
        x"940E",
        x"047B",
        x"E385",
        x"958A",
        x"F7F1",
        x"E082",
        x"E090",
        x"940E",
        x"0494",
        x"9508",
        x"B392",
        x"7C90",
        x"BB92",
        x"B392",
        x"2B98",
        x"BB92",
        x"E085",
        x"958A",
        x"F7F1",
        x"0000",
        x"B181",
        x"9A90",
        x"E095",
        x"959A",
        x"F7F1",
        x"0000",
        x"B121",
        x"E090",
        x"2B92",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2FC6",
        x"2FD7",
        x"161C",
        x"061D",
        x"F464",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E084",
        x"E090",
        x"940E",
        x"047B",
        x"9516",
        x"9507",
        x"9721",
        x"CFF1",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC6",
        x"2FD7",
        x"2EE4",
        x"2EF5",
        x"2F02",
        x"2F13",
        x"E160",
        x"E070",
        x"940E",
        x"04D1",
        x"E160",
        x"E070",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"04D1",
        x"E06A",
        x"E070",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"04D1",
        x"E064",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"04D1",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"14F0",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"E0C8",
        x"E0D0",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E08C",
        x"E090",
        x"940E",
        x"047B",
        x"9516",
        x"9507",
        x"9721",
        x"9720",
        x"F799",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"E1C0",
        x"E0D0",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E08C",
        x"E090",
        x"940E",
        x"047B",
        x"9516",
        x"9507",
        x"9721",
        x"9720",
        x"F799",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"93CF",
        x"93DF",
        x"E02C",
        x"E033",
        x"933F",
        x"932F",
        x"E22A",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"9180",
        x"030C",
        x"9190",
        x"030D",
        x"940E",
        x"052E",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E0CA",
        x"E0D0",
        x"9180",
        x"030C",
        x"9190",
        x"030D",
        x"940E",
        x"11FA",
        x"9390",
        x"030D",
        x"9380",
        x"030C",
        x"9721",
        x"9720",
        x"F799",
        x"91DF",
        x"91CF",
        x"9508",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2D",
        x"4F3F",
        x"933F",
        x"932F",
        x"E227",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"818B",
        x"819C",
        x"940E",
        x"052E",
        x"804B",
        x"805C",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2C81",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"2C61",
        x"2C71",
        x"8189",
        x"819A",
        x"E0A0",
        x"E0B0",
        x"2D7B",
        x"2D6A",
        x"2D59",
        x"2D48",
        x"0D44",
        x"1D55",
        x"1D66",
        x"1D77",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F154",
        x"940E",
        x"04AF",
        x"E028",
        x"E030",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"0F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"2EC8",
        x"2ED9",
        x"E0E1",
        x"22CE",
        x"24DD",
        x"2CE1",
        x"2CF1",
        x"2AC4",
        x"2AD5",
        x"2AE6",
        x"2AF7",
        x"9596",
        x"9587",
        x"FEE0",
        x"C004",
        x"E24D",
        x"26C4",
        x"24EE",
        x"24FF",
        x"5021",
        x"0931",
        x"1521",
        x"0531",
        x"F701",
        x"EF8F",
        x"1A88",
        x"0A98",
        x"0AA8",
        x"0AB8",
        x"CFC5",
        x"92FF",
        x"92EF",
        x"92DF",
        x"92CF",
        x"E58A",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"9508",
        x"E060",
        x"E070",
        x"E183",
        x"E090",
        x"940E",
        x"047B",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2D",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2B",
        x"4F3F",
        x"933F",
        x"932F",
        x"E224",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"818A",
        x"938F",
        x"8189",
        x"938F",
        x"818C",
        x"938F",
        x"818B",
        x"938F",
        x"818E",
        x"938F",
        x"818D",
        x"938F",
        x"E685",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"8189",
        x"819A",
        x"940E",
        x"0514",
        x"818D",
        x"819E",
        x"940E",
        x"052E",
        x"808D",
        x"809E",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"2CA1",
        x"2CB1",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"0D48",
        x"1D59",
        x"1D6A",
        x"1D7B",
        x"EF9F",
        x"1AC9",
        x"0AD9",
        x"0AE9",
        x"0AF9",
        x"818B",
        x"819C",
        x"E0A0",
        x"E0B0",
        x"1784",
        x"0795",
        x"07A6",
        x"07B7",
        x"F01C",
        x"940E",
        x"0610",
        x"CFE7",
        x"9626",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"E060",
        x"E070",
        x"E184",
        x"E090",
        x"940E",
        x"047B",
        x"E385",
        x"958A",
        x"F7F1",
        x"E082",
        x"E090",
        x"940E",
        x"0494",
        x"9508",
        x"E060",
        x"E070",
        x"E185",
        x"E090",
        x"940E",
        x"047B",
        x"E385",
        x"958A",
        x"F7F1",
        x"E082",
        x"E090",
        x"940E",
        x"0494",
        x"9508",
        x"E060",
        x"E070",
        x"E186",
        x"E090",
        x"940E",
        x"047B",
        x"9508",
        x"E060",
        x"E070",
        x"E187",
        x"E090",
        x"940E",
        x"047B",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"052E",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"11FA",
        x"91DF",
        x"91CF",
        x"9508",
        x"E2A2",
        x"E0B0",
        x"EDE2",
        x"E0F6",
        x"940C",
        x"14C8",
        x"A37A",
        x"A369",
        x"E02C",
        x"E033",
        x"933F",
        x"932F",
        x"E22A",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"9180",
        x"030C",
        x"9190",
        x"030D",
        x"940E",
        x"052E",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2CE1",
        x"2CF1",
        x"2EAC",
        x"2EBD",
        x"E221",
        x"0EA2",
        x"1CB1",
        x"E102",
        x"E011",
        x"EFAC",
        x"2E2A",
        x"E0A3",
        x"2E3A",
        x"2EC0",
        x"2ED1",
        x"EFBA",
        x"2E4B",
        x"E0B3",
        x"2E5B",
        x"EF87",
        x"2E68",
        x"E083",
        x"2E78",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2E88",
        x"2E99",
        x"A1E9",
        x"A1FA",
        x"9509",
        x"2DA8",
        x"2DB9",
        x"938D",
        x"939D",
        x"2E8A",
        x"2E9B",
        x"15AA",
        x"05BB",
        x"F7A1",
        x"9180",
        x"030C",
        x"9190",
        x"030D",
        x"0D8E",
        x"1D9F",
        x"939F",
        x"938F",
        x"E0A2",
        x"E0B4",
        x"93BF",
        x"93AF",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2E88",
        x"2E99",
        x"2DA8",
        x"2DB9",
        x"918C",
        x"9611",
        x"919C",
        x"E0B2",
        x"0E8B",
        x"1C91",
        x"939F",
        x"938F",
        x"923F",
        x"922F",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"148A",
        x"049B",
        x"F739",
        x"925F",
        x"924F",
        x"92DF",
        x"92CF",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2FEC",
        x"2FFD",
        x"9631",
        x"2E8E",
        x"2E9F",
        x"2DA8",
        x"2DB9",
        x"918D",
        x"919D",
        x"2E8A",
        x"2E9B",
        x"2F48",
        x"2F59",
        x"5240",
        x"0951",
        x"354F",
        x"0551",
        x"F010",
        x"E28E",
        x"E090",
        x"939F",
        x"938F",
        x"927F",
        x"926F",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"148A",
        x"049B",
        x"F701",
        x"EFA5",
        x"E0B3",
        x"93BF",
        x"93AF",
        x"92DF",
        x"92CF",
        x"940E",
        x"1579",
        x"E1F0",
        x"0EEF",
        x"1CF1",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"14E1",
        x"E021",
        x"06F2",
        x"F009",
        x"CF78",
        x"9180",
        x"030C",
        x"9190",
        x"030D",
        x"9593",
        x"9390",
        x"030D",
        x"9380",
        x"030C",
        x"96A2",
        x"E1E2",
        x"940C",
        x"14E4",
        x"EA6F",
        x"E074",
        x"940E",
        x"06CC",
        x"9508",
        x"E0A8",
        x"E0B0",
        x"EAE3",
        x"E0F7",
        x"940C",
        x"14D6",
        x"2F06",
        x"2F17",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2B",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F29",
        x"4F3F",
        x"933F",
        x"932F",
        x"E22D",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"818E",
        x"938F",
        x"818D",
        x"938F",
        x"8588",
        x"938F",
        x"818F",
        x"938F",
        x"EE84",
        x"E093",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"818D",
        x"819E",
        x"940E",
        x"0514",
        x"818F",
        x"8598",
        x"940E",
        x"052E",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"5041",
        x"0951",
        x"0961",
        x"0971",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"1618",
        x"0619",
        x"061A",
        x"061B",
        x"F424",
        x"2FE0",
        x"2FF1",
        x"9509",
        x"CFE7",
        x"9628",
        x"E0E4",
        x"940C",
        x"14F2",
        x"E86D",
        x"E074",
        x"940E",
        x"079D",
        x"9508",
        x"E0A6",
        x"E0B0",
        x"E0EE",
        x"E0F8",
        x"940C",
        x"14CE",
        x"2F06",
        x"2F17",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2B",
        x"4F3F",
        x"933F",
        x"932F",
        x"E320",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"818D",
        x"819E",
        x"940E",
        x"052E",
        x"2FE0",
        x"2FF1",
        x"9509",
        x"2EA8",
        x"2EB9",
        x"92BF",
        x"938F",
        x"818E",
        x"938F",
        x"818D",
        x"938F",
        x"ED83",
        x"E093",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"EB94",
        x"2EE9",
        x"E093",
        x"2EF9",
        x"E122",
        x"2EC2",
        x"E021",
        x"2ED2",
        x"8149",
        x"815A",
        x"816B",
        x"817C",
        x"2FB7",
        x"2FA6",
        x"2F95",
        x"2F84",
        x"9701",
        x"09A1",
        x"09B1",
        x"8389",
        x"839A",
        x"83AB",
        x"83BC",
        x"3042",
        x"0551",
        x"0561",
        x"0571",
        x"F0D4",
        x"2FE0",
        x"2FF1",
        x"9509",
        x"2E88",
        x"2E99",
        x"158A",
        x"059B",
        x"F079",
        x"92BF",
        x"92AF",
        x"929F",
        x"938F",
        x"92FF",
        x"92EF",
        x"92DF",
        x"92CF",
        x"940E",
        x"1579",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2CA8",
        x"2CB9",
        x"CFD2",
        x"9626",
        x"E0EC",
        x"940C",
        x"14EA",
        x"EA61",
        x"E074",
        x"940E",
        x"0808",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2F86",
        x"2F97",
        x"940E",
        x"0494",
        x"2FC8",
        x"2FD9",
        x"2F80",
        x"2F91",
        x"940E",
        x"04BD",
        x"2F08",
        x"2F19",
        x"2F8C",
        x"2F9D",
        x"E0A0",
        x"E0B0",
        x"2777",
        x"2766",
        x"E020",
        x"E030",
        x"2B60",
        x"2B71",
        x"2B82",
        x"2B93",
        x"E420",
        x"E432",
        x"E04F",
        x"E050",
        x"940E",
        x"14A1",
        x"939F",
        x"938F",
        x"937F",
        x"936F",
        x"935F",
        x"934F",
        x"933F",
        x"932F",
        x"EA86",
        x"E093",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"B78D",
        x"B79E",
        x"960C",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"EDE2",
        x"E0F8",
        x"940C",
        x"14D0",
        x"2EE8",
        x"2EF9",
        x"E9C0",
        x"E0D0",
        x"E081",
        x"E090",
        x"EA50",
        x"2EC5",
        x"E053",
        x"2ED5",
        x"E102",
        x"E011",
        x"EA63",
        x"2EA6",
        x"E063",
        x"2EB6",
        x"FEE0",
        x"C01E",
        x"2B89",
        x"F451",
        x"92BF",
        x"92AF",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"8189",
        x"938F",
        x"8188",
        x"938F",
        x"92DF",
        x"92CF",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E080",
        x"E090",
        x"94F6",
        x"94E7",
        x"9622",
        x"E020",
        x"3AC4",
        x"07D2",
        x"F6C9",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"14EC",
        x"3180",
        x"0591",
        x"F4D8",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"59E0",
        x"4FFF",
        x"8181",
        x"938F",
        x"8180",
        x"938F",
        x"E984",
        x"E093",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"E883",
        x"E093",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E4E1",
        x"E0F9",
        x"940C",
        x"14C8",
        x"9180",
        x"030E",
        x"9190",
        x"030F",
        x"2B89",
        x"F409",
        x"C069",
        x"E4E4",
        x"2E6E",
        x"E0E3",
        x"2E7E",
        x"E5F4",
        x"2E4F",
        x"E0F3",
        x"2E5F",
        x"E6A4",
        x"2EEA",
        x"E0A3",
        x"2EFA",
        x"E3B0",
        x"2ECB",
        x"E0B3",
        x"2EDB",
        x"E000",
        x"E010",
        x"E4C5",
        x"2E2C",
        x"E0C1",
        x"2E3C",
        x"E1C2",
        x"E0D1",
        x"E482",
        x"2EA8",
        x"E081",
        x"2EB8",
        x"E39F",
        x"2E89",
        x"E091",
        x"2E99",
        x"9180",
        x"030E",
        x"9190",
        x"030F",
        x"1708",
        x"0719",
        x"F00C",
        x"C04F",
        x"2DE6",
        x"2DF7",
        x"8120",
        x"8131",
        x"E0F2",
        x"0E6F",
        x"1C71",
        x"2DE4",
        x"2DF5",
        x"8180",
        x"8191",
        x"E0F2",
        x"0E4F",
        x"1C51",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"923F",
        x"922F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"2DEE",
        x"2DFF",
        x"9181",
        x"9191",
        x"2EEE",
        x"2EFF",
        x"940E",
        x"08CC",
        x"92BF",
        x"92AF",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"2DEC",
        x"2DFD",
        x"9181",
        x"9191",
        x"2ECE",
        x"2EDF",
        x"940E",
        x"090E",
        x"929F",
        x"928F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"5F0F",
        x"4F1F",
        x"B78D",
        x"B79E",
        x"9642",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"CFB7",
        x"E28B",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E1E2",
        x"940C",
        x"14E4",
        x"E0A0",
        x"E0B0",
        x"ECEA",
        x"E0F9",
        x"940C",
        x"14CE",
        x"E086",
        x"E090",
        x"940E",
        x"04BD",
        x"2EC8",
        x"2ED9",
        x"E088",
        x"E090",
        x"940E",
        x"04BD",
        x"2EB8",
        x"2EA9",
        x"E08A",
        x"E090",
        x"940E",
        x"0494",
        x"2E98",
        x"2E89",
        x"E08B",
        x"E090",
        x"940E",
        x"0494",
        x"2EE8",
        x"2EF9",
        x"E021",
        x"22E2",
        x"24FF",
        x"E001",
        x"E010",
        x"C002",
        x"0F00",
        x"1F11",
        x"958A",
        x"F7E2",
        x"2F80",
        x"2F91",
        x"7A8A",
        x"7092",
        x"2B89",
        x"F031",
        x"E06E",
        x"E070",
        x"E08C",
        x"E090",
        x"940E",
        x"0889",
        x"2F80",
        x"2F91",
        x"940E",
        x"08CC",
        x"92DF",
        x"92CF",
        x"E726",
        x"E033",
        x"933F",
        x"932F",
        x"E1C2",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2300",
        x"F181",
        x"2F80",
        x"2F91",
        x"7C8C",
        x"2799",
        x"2B89",
        x"F039",
        x"E62D",
        x"E033",
        x"933F",
        x"932F",
        x"93DF",
        x"93CF",
        x"C006",
        x"E624",
        x"E033",
        x"933F",
        x"932F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"E526",
        x"E033",
        x"933F",
        x"932F",
        x"E122",
        x"E031",
        x"933F",
        x"932F",
        x"940E",
        x"1579",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C00C",
        x"E524",
        x"E033",
        x"933F",
        x"932F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"7505",
        x"2711",
        x"1501",
        x"0511",
        x"F051",
        x"E06E",
        x"E070",
        x"E08C",
        x"E090",
        x"940E",
        x"0889",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"06BF",
        x"2D8E",
        x"2D9F",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"14EA",
        x"E080",
        x"E090",
        x"940E",
        x"04BD",
        x"9390",
        x"030D",
        x"9380",
        x"030C",
        x"E063",
        x"E070",
        x"E084",
        x"E090",
        x"940E",
        x"0889",
        x"9180",
        x"030C",
        x"9190",
        x"030D",
        x"940E",
        x"06BF",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"E620",
        x"E030",
        x"933F",
        x"932F",
        x"E323",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"9180",
        x"0060",
        x"9190",
        x"0061",
        x"91A0",
        x"0062",
        x"91B0",
        x"0063",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"1618",
        x"0619",
        x"061A",
        x"061B",
        x"F07C",
        x"EA88",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C06C",
        x"93BF",
        x"93AF",
        x"939F",
        x"938F",
        x"E88D",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"9080",
        x"0340",
        x"9090",
        x"0341",
        x"90A0",
        x"0342",
        x"90B0",
        x"0343",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"24CC",
        x"94C3",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"9180",
        x"0060",
        x"9190",
        x"0061",
        x"91A0",
        x"0062",
        x"91B0",
        x"0063",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F1E4",
        x"E060",
        x"E070",
        x"E088",
        x"E090",
        x"940E",
        x"047B",
        x"9180",
        x"0060",
        x"9190",
        x"0061",
        x"91A0",
        x"0062",
        x"91B0",
        x"0063",
        x"16C8",
        x"06D9",
        x"06EA",
        x"06FB",
        x"F0B1",
        x"9180",
        x"0340",
        x"9190",
        x"0341",
        x"91A0",
        x"0342",
        x"91B0",
        x"0343",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F0B9",
        x"E091",
        x"1A89",
        x"0891",
        x"08A1",
        x"08B1",
        x"1481",
        x"0491",
        x"04A1",
        x"04B1",
        x"F469",
        x"E385",
        x"958A",
        x"F7F1",
        x"940E",
        x"0A62",
        x"9080",
        x"0340",
        x"9090",
        x"0341",
        x"90A0",
        x"0342",
        x"90B0",
        x"0343",
        x"EF9F",
        x"1AC9",
        x"0AD9",
        x"0AE9",
        x"0AF9",
        x"CFB7",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"93CF",
        x"93DF",
        x"E78E",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E0C2",
        x"E0D0",
        x"E061",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"047B",
        x"EC86",
        x"E090",
        x"9701",
        x"F7F1",
        x"E060",
        x"E070",
        x"E088",
        x"E090",
        x"940E",
        x"047B",
        x"EC86",
        x"E090",
        x"9701",
        x"F7F1",
        x"E060",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"047B",
        x"EC86",
        x"E090",
        x"9701",
        x"F7F1",
        x"9721",
        x"9720",
        x"F6F9",
        x"940E",
        x"0A62",
        x"91DF",
        x"91CF",
        x"9508",
        x"93CF",
        x"93DF",
        x"E387",
        x"E091",
        x"939F",
        x"938F",
        x"E38C",
        x"E091",
        x"939F",
        x"938F",
        x"E381",
        x"E093",
        x"939F",
        x"938F",
        x"E1C2",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"E484",
        x"E091",
        x"939F",
        x"938F",
        x"E580",
        x"E091",
        x"939F",
        x"938F",
        x"E18B",
        x"E093",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"921F",
        x"E088",
        x"938F",
        x"EF87",
        x"E092",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"B78D",
        x"B79E",
        x"9646",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"940E",
        x"0B5A",
        x"ED88",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"EDC0",
        x"E0D0",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"ED30",
        x"2EE3",
        x"E031",
        x"2EF3",
        x"E102",
        x"E011",
        x"8188",
        x"8199",
        x"9622",
        x"939F",
        x"938F",
        x"92FF",
        x"92EF",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E080",
        x"3FCC",
        x"07D8",
        x"F759",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"14F0",
        x"E0A2",
        x"E0B0",
        x"EDE2",
        x"E0FB",
        x"940C",
        x"14D8",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E22A",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"9140",
        x"030E",
        x"9150",
        x"030F",
        x"8129",
        x"813A",
        x"E5E4",
        x"E0F3",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E080",
        x"E090",
        x"1784",
        x"0795",
        x"F454",
        x"9161",
        x"9171",
        x"1762",
        x"0773",
        x"F419",
        x"839A",
        x"8389",
        x"C002",
        x"9601",
        x"CFF3",
        x"8129",
        x"813A",
        x"1724",
        x"0735",
        x"F0AC",
        x"933F",
        x"932F",
        x"ED85",
        x"E092",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"EF8F",
        x"EF9F",
        x"C002",
        x"2F82",
        x"2F93",
        x"9622",
        x"E0E2",
        x"940C",
        x"14F4",
        x"E0A0",
        x"E0B0",
        x"E2E7",
        x"E0FC",
        x"940C",
        x"14D0",
        x"940E",
        x"0BCC",
        x"2FC8",
        x"2FD9",
        x"FD97",
        x"C085",
        x"E281",
        x"E091",
        x"939F",
        x"938F",
        x"E142",
        x"2EE4",
        x"E041",
        x"2EF4",
        x"92FF",
        x"92EF",
        x"940E",
        x"1579",
        x"2F0C",
        x"2F1D",
        x"0F00",
        x"1F11",
        x"2F20",
        x"2F31",
        x"592C",
        x"4F3C",
        x"2EA2",
        x"2EB3",
        x"2FE2",
        x"2FF3",
        x"8180",
        x"8191",
        x"940E",
        x"08CC",
        x"2F20",
        x"2F31",
        x"5A2C",
        x"4F3C",
        x"2EC2",
        x"2ED3",
        x"2FE2",
        x"2FF3",
        x"8181",
        x"938F",
        x"8180",
        x"938F",
        x"E187",
        x"E091",
        x"939F",
        x"938F",
        x"92FF",
        x"92EF",
        x"940E",
        x"1579",
        x"9180",
        x"030E",
        x"9190",
        x"030F",
        x"2F60",
        x"2F71",
        x"5B6C",
        x"4F7C",
        x"5D00",
        x"4F1C",
        x"B72D",
        x"B73E",
        x"5F26",
        x"4F3F",
        x"B60F",
        x"94F8",
        x"BF3E",
        x"BE0F",
        x"BF2D",
        x"E040",
        x"E050",
        x"E020",
        x"E030",
        x"5F2E",
        x"4F3F",
        x"17C8",
        x"07D9",
        x"F5A4",
        x"9621",
        x"2DEC",
        x"2DFD",
        x"0FE2",
        x"1FF3",
        x"81A0",
        x"81B1",
        x"2DEC",
        x"2DFD",
        x"0FE4",
        x"1FF5",
        x"83B1",
        x"83A0",
        x"2FE6",
        x"2FF7",
        x"0FE2",
        x"1FF3",
        x"81A0",
        x"81B1",
        x"2FE6",
        x"2FF7",
        x"0FE4",
        x"1FF5",
        x"83B1",
        x"83A0",
        x"2DEA",
        x"2DFB",
        x"0FE2",
        x"1FF3",
        x"81A0",
        x"81B1",
        x"2DEA",
        x"2DFB",
        x"0FE4",
        x"1FF5",
        x"83B1",
        x"83A0",
        x"2FE0",
        x"2FF1",
        x"0FE2",
        x"1FF3",
        x"81A0",
        x"81B1",
        x"2FE0",
        x"2FF1",
        x"0FE4",
        x"1FF5",
        x"83B1",
        x"83A0",
        x"5F4E",
        x"4F5F",
        x"CFC7",
        x"9701",
        x"9390",
        x"030F",
        x"9380",
        x"030E",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"14EC",
        x"E0A2",
        x"E0B0",
        x"EBED",
        x"E0FC",
        x"940C",
        x"14D4",
        x"2EF8",
        x"2EE9",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"940E",
        x"0BCC",
        x"2F08",
        x"2F19",
        x"FF97",
        x"C039",
        x"E087",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"821A",
        x"8219",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"EF0A",
        x"E010",
        x"E1E2",
        x"2EEE",
        x"E0E1",
        x"2EFE",
        x"8189",
        x"819A",
        x"3180",
        x"0591",
        x"F00C",
        x"C04D",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"59E0",
        x"4FFF",
        x"8121",
        x"932F",
        x"8120",
        x"932F",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"92FF",
        x"92EF",
        x"940E",
        x"1579",
        x"8189",
        x"819A",
        x"9601",
        x"839A",
        x"8389",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"CFDD",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E529",
        x"E031",
        x"933F",
        x"932F",
        x"92EF",
        x"92FF",
        x"940E",
        x"1598",
        x"8189",
        x"819A",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"3180",
        x"0591",
        x"F448",
        x"2FE0",
        x"2FF1",
        x"0FEE",
        x"1FFF",
        x"5DE0",
        x"4FFC",
        x"8391",
        x"8380",
        x"C00E",
        x"EC87",
        x"E090",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9622",
        x"E0E6",
        x"940C",
        x"14F0",
        x"E061",
        x"E070",
        x"2B89",
        x"F411",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"047B",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"E4E7",
        x"E0FD",
        x"940C",
        x"14CC",
        x"821A",
        x"8219",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E626",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"E060",
        x"E070",
        x"E082",
        x"E090",
        x"940E",
        x"047B",
        x"E3F0",
        x"2E6F",
        x"E0F3",
        x"2E7F",
        x"E6A4",
        x"2EAA",
        x"E0A3",
        x"2EBA",
        x"E4B4",
        x"2ECB",
        x"E0B3",
        x"2EDB",
        x"E514",
        x"2E81",
        x"E013",
        x"2E91",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2CE1",
        x"2CF1",
        x"9100",
        x"030E",
        x"9110",
        x"030F",
        x"16E0",
        x"06F1",
        x"F4F4",
        x"2DE6",
        x"2DF7",
        x"9121",
        x"9131",
        x"2E6E",
        x"2E7F",
        x"2DEA",
        x"2DFB",
        x"9141",
        x"9151",
        x"2EAE",
        x"2EBF",
        x"2DEC",
        x"2DFD",
        x"9161",
        x"9171",
        x"2ECE",
        x"2EDF",
        x"2DE8",
        x"2DF9",
        x"9181",
        x"9191",
        x"2E8E",
        x"2E9F",
        x"940E",
        x"04ED",
        x"EFFF",
        x"1AEF",
        x"0AFF",
        x"CFDB",
        x"3008",
        x"0511",
        x"F46C",
        x"E020",
        x"E030",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"04ED",
        x"5F0F",
        x"4F1F",
        x"CFF0",
        x"E060",
        x"E070",
        x"E088",
        x"E090",
        x"940E",
        x"047B",
        x"E061",
        x"E070",
        x"E082",
        x"E090",
        x"940E",
        x"047B",
        x"E080",
        x"E090",
        x"940E",
        x"0D36",
        x"8189",
        x"819A",
        x"2B89",
        x"F0F9",
        x"EB88",
        x"E090",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"E061",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"047B",
        x"E88C",
        x"E091",
        x"9701",
        x"F7F1",
        x"0000",
        x"E060",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"047B",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"EA83",
        x"E090",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E001",
        x"E010",
        x"B2F0",
        x"FEF7",
        x"C00A",
        x"940E",
        x"09C4",
        x"2F08",
        x"2F19",
        x"E060",
        x"E070",
        x"E089",
        x"E090",
        x"940E",
        x"047B",
        x"FEF6",
        x"C002",
        x"E000",
        x"E010",
        x"940E",
        x"1468",
        x"2388",
        x"F031",
        x"940E",
        x"1462",
        x"308D",
        x"F411",
        x"E000",
        x"E010",
        x"E395",
        x"959A",
        x"F7F1",
        x"1501",
        x"0511",
        x"F6F9",
        x"E986",
        x"E090",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"E081",
        x"E090",
        x"940E",
        x"0D36",
        x"E060",
        x"E070",
        x"E082",
        x"E090",
        x"940E",
        x"047B",
        x"940E",
        x"0A62",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9622",
        x"E0EE",
        x"940C",
        x"14E8",
        x"9360",
        x"0340",
        x"9370",
        x"0341",
        x"9380",
        x"0342",
        x"9390",
        x"0343",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F0B9",
        x"939F",
        x"938F",
        x"937F",
        x"936F",
        x"E98F",
        x"E092",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"9508",
        x"E88D",
        x"E092",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"E6E5",
        x"E0FE",
        x"940C",
        x"14D8",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"E323",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"8169",
        x"817A",
        x"818B",
        x"819C",
        x"940E",
        x"0E2C",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"9624",
        x"E0E2",
        x"940C",
        x"14F4",
        x"E0A0",
        x"E0B0",
        x"E8E9",
        x"E0FE",
        x"940C",
        x"14D0",
        x"2EA8",
        x"2EB9",
        x"2FC6",
        x"2FD7",
        x"2EE4",
        x"2EF5",
        x"2EC2",
        x"2ED3",
        x"2F82",
        x"2F93",
        x"940E",
        x"08CC",
        x"93DF",
        x"93CF",
        x"E78F",
        x"E092",
        x"939F",
        x"938F",
        x"E122",
        x"E031",
        x"933F",
        x"932F",
        x"940E",
        x"1579",
        x"2DEA",
        x"2DFB",
        x"0FEE",
        x"1FFF",
        x"2FAE",
        x"2FBF",
        x"5AAC",
        x"4FBC",
        x"21CE",
        x"21DF",
        x"93CD",
        x"93DC",
        x"2FAE",
        x"2FBF",
        x"5BAC",
        x"4FBC",
        x"92ED",
        x"92FC",
        x"2FAE",
        x"2FBF",
        x"59AC",
        x"4FBC",
        x"92CD",
        x"92DC",
        x"5DE0",
        x"4FFC",
        x"8311",
        x"8300",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"14EC",
        x"E0A6",
        x"E0B0",
        x"ECEE",
        x"E0FE",
        x"940C",
        x"14CC",
        x"2EE6",
        x"2EF7",
        x"EF2F",
        x"EF3F",
        x"833C",
        x"832B",
        x"833A",
        x"8329",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2D",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2B",
        x"4F3F",
        x"933F",
        x"932F",
        x"E224",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"9120",
        x"030E",
        x"9130",
        x"030F",
        x"816D",
        x"817E",
        x"E5E4",
        x"E0F3",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"E080",
        x"E090",
        x"1782",
        x"0793",
        x"F5AC",
        x"9141",
        x"9151",
        x"1746",
        x"0757",
        x"F571",
        x"2F48",
        x"2F59",
        x"0F44",
        x"1F55",
        x"2FE4",
        x"2FF5",
        x"59EC",
        x"4FFC",
        x"8120",
        x"8131",
        x"2FE2",
        x"2FF3",
        x"21EE",
        x"21FF",
        x"2BEF",
        x"F059",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"08CC",
        x"818E",
        x"938F",
        x"818D",
        x"938F",
        x"E689",
        x"E092",
        x"C01D",
        x"81E9",
        x"81FA",
        x"9631",
        x"F441",
        x"2FE4",
        x"2FF5",
        x"5DE0",
        x"4FFC",
        x"8140",
        x"8151",
        x"835A",
        x"8349",
        x"8109",
        x"811A",
        x"292E",
        x"293F",
        x"814B",
        x"815C",
        x"C0A4",
        x"9601",
        x"CFC8",
        x"3028",
        x"0531",
        x"F4A1",
        x"921F",
        x"E088",
        x"938F",
        x"E485",
        x"E092",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C08D",
        x"2F82",
        x"2F93",
        x"9601",
        x"9390",
        x"030F",
        x"9380",
        x"030E",
        x"8189",
        x"819A",
        x"9601",
        x"F421",
        x"E08F",
        x"E090",
        x"839A",
        x"8389",
        x"2E62",
        x"2E73",
        x"E011",
        x"1A61",
        x"0871",
        x"2F82",
        x"2F93",
        x"0F88",
        x"1F99",
        x"2F28",
        x"2F39",
        x"5A2C",
        x"4F3C",
        x"2F48",
        x"2F59",
        x"5B4C",
        x"4F5C",
        x"2E84",
        x"2E95",
        x"2FA8",
        x"2FB9",
        x"59AC",
        x"4FBC",
        x"2EAA",
        x"2EBB",
        x"5D80",
        x"4F9C",
        x"E0E2",
        x"E0F0",
        x"E040",
        x"E050",
        x"C04A",
        x"9732",
        x"5042",
        x"0951",
        x"2F02",
        x"2F13",
        x"0F04",
        x"1F15",
        x"2FA0",
        x"2FB1",
        x"910D",
        x"911C",
        x"1706",
        x"0717",
        x"F408",
        x"C044",
        x"2EC2",
        x"2ED3",
        x"0ECE",
        x"1EDF",
        x"2DAC",
        x"2DBD",
        x"930D",
        x"931C",
        x"2D08",
        x"2D19",
        x"0F04",
        x"1F15",
        x"2FA0",
        x"2FB1",
        x"90CD",
        x"90DC",
        x"2D08",
        x"2D19",
        x"0F0E",
        x"1F1F",
        x"2FA0",
        x"2FB1",
        x"92CD",
        x"92DC",
        x"2D0A",
        x"2D1B",
        x"0F04",
        x"1F15",
        x"2FA0",
        x"2FB1",
        x"90CD",
        x"90DC",
        x"2D0A",
        x"2D1B",
        x"0F0E",
        x"1F1F",
        x"2FA0",
        x"2FB1",
        x"92CD",
        x"92DC",
        x"2F08",
        x"2F19",
        x"0F04",
        x"1F15",
        x"2FA0",
        x"2FB1",
        x"90CD",
        x"90DC",
        x"2F08",
        x"2F19",
        x"0F0E",
        x"1F1F",
        x"2FA0",
        x"2FB1",
        x"92CD",
        x"92DC",
        x"E0B1",
        x"1A6B",
        x"0871",
        x"EF1F",
        x"1661",
        x"0671",
        x"F084",
        x"EFBF",
        x"166B",
        x"067B",
        x"F009",
        x"CFAD",
        x"8109",
        x"811A",
        x"814B",
        x"815C",
        x"2D2E",
        x"2D3F",
        x"2D86",
        x"2D97",
        x"9601",
        x"940E",
        x"0E83",
        x"9626",
        x"E0EE",
        x"940C",
        x"14E8",
        x"E060",
        x"E071",
        x"940E",
        x"0EC8",
        x"9508",
        x"E060",
        x"E072",
        x"940E",
        x"0EC8",
        x"9508",
        x"E061",
        x"E070",
        x"940E",
        x"0EC8",
        x"9508",
        x"E062",
        x"E070",
        x"940E",
        x"0EC8",
        x"9508",
        x"E064",
        x"E070",
        x"940E",
        x"0EC8",
        x"9508",
        x"E068",
        x"E070",
        x"940E",
        x"0EC8",
        x"9508",
        x"3F6F",
        x"EF2F",
        x"0772",
        x"F419",
        x"FF80",
        x"C026",
        x"C028",
        x"3F6E",
        x"EF4F",
        x"0774",
        x"F419",
        x"FF80",
        x"C022",
        x"C01E",
        x"3F6D",
        x"EF2F",
        x"0772",
        x"F429",
        x"2F28",
        x"2F39",
        x"EC43",
        x"2724",
        x"C008",
        x"3F6C",
        x"EF2F",
        x"0772",
        x"F441",
        x"2F28",
        x"2F39",
        x"E34C",
        x"2724",
        x"2F89",
        x"2799",
        x"2782",
        x"9508",
        x"FF77",
        x"C003",
        x"940E",
        x"1559",
        x"C002",
        x"2F86",
        x"2F97",
        x"2799",
        x"9508",
        x"EA8A",
        x"E090",
        x"9508",
        x"E585",
        x"E090",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E3E5",
        x"E1F0",
        x"940C",
        x"14C8",
        x"2F08",
        x"2F19",
        x"2E46",
        x"2E57",
        x"2FC4",
        x"2FD5",
        x"2F84",
        x"2F95",
        x"940E",
        x"155E",
        x"2EC0",
        x"2ED1",
        x"2CE1",
        x"2CF1",
        x"2C81",
        x"2C91",
        x"2CA1",
        x"2CB1",
        x"2C61",
        x"2C71",
        x"2DBB",
        x"2DAA",
        x"2D99",
        x"2D88",
        x"0D8C",
        x"1D9D",
        x"1DAE",
        x"1DBF",
        x"1648",
        x"0659",
        x"066A",
        x"067B",
        x"F0C4",
        x"2E20",
        x"2E31",
        x"0C28",
        x"1C39",
        x"2F6C",
        x"2F7D",
        x"2D82",
        x"2D93",
        x"940E",
        x"0FFD",
        x"940E",
        x"0514",
        x"2D82",
        x"2D93",
        x"940E",
        x"052E",
        x"940E",
        x"0610",
        x"EF8F",
        x"1A88",
        x"0A98",
        x"0AA8",
        x"0AB8",
        x"CFDB",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"155E",
        x"2F80",
        x"2F91",
        x"940E",
        x"052E",
        x"2C21",
        x"2C31",
        x"E108",
        x"E012",
        x"E162",
        x"2EA6",
        x"E061",
        x"2EB6",
        x"144C",
        x"045D",
        x"046E",
        x"047F",
        x"F164",
        x"940E",
        x"04AF",
        x"2E88",
        x"2E99",
        x"2F6C",
        x"2F7D",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"0FFD",
        x"1588",
        x"0599",
        x"F0C9",
        x"929F",
        x"928F",
        x"939F",
        x"938F",
        x"92FF",
        x"92EF",
        x"92DF",
        x"92CF",
        x"931F",
        x"930F",
        x"92BF",
        x"92AF",
        x"940E",
        x"1579",
        x"EF9F",
        x"1A29",
        x"0A39",
        x"B78D",
        x"B79E",
        x"960C",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"EF9F",
        x"1AC9",
        x"0AD9",
        x"0AE9",
        x"0AF9",
        x"CFCF",
        x"2788",
        x"2799",
        x"1B8C",
        x"0B9D",
        x"FD97",
        x"C006",
        x"3086",
        x"0591",
        x"F02C",
        x"E085",
        x"E090",
        x"C002",
        x"E080",
        x"E090",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"59EC",
        x"4FFF",
        x"8181",
        x"938F",
        x"8180",
        x"938F",
        x"E088",
        x"E092",
        x"939F",
        x"938F",
        x"E102",
        x"E011",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"FDD7",
        x"C010",
        x"93DF",
        x"93CF",
        x"E082",
        x"E092",
        x"939F",
        x"938F",
        x"931F",
        x"930F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"1421",
        x"0431",
        x"F099",
        x"923F",
        x"922F",
        x"EE8D",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C00E",
        x"EE83",
        x"E091",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E1E2",
        x"940C",
        x"14E4",
        x"E0A6",
        x"E0B0",
        x"E1E8",
        x"E1F1",
        x"940C",
        x"14D6",
        x"E92C",
        x"EF3F",
        x"833A",
        x"8329",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2D",
        x"4F3F",
        x"933F",
        x"932F",
        x"2F2C",
        x"2F3D",
        x"5F2B",
        x"4F3F",
        x"933F",
        x"932F",
        x"E620",
        x"E031",
        x"933F",
        x"932F",
        x"939F",
        x"938F",
        x"940E",
        x"1598",
        x"8149",
        x"815A",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"816B",
        x"817C",
        x"818D",
        x"819E",
        x"394C",
        x"EF2F",
        x"0752",
        x"F529",
        x"E545",
        x"E050",
        x"940E",
        x"102F",
        x"816B",
        x"817C",
        x"EA4A",
        x"E050",
        x"818D",
        x"819E",
        x"940E",
        x"102F",
        x"816B",
        x"817C",
        x"EF4F",
        x"E050",
        x"818D",
        x"819E",
        x"940E",
        x"102F",
        x"E000",
        x"E010",
        x"816B",
        x"817C",
        x"2F40",
        x"2F51",
        x"818D",
        x"819E",
        x"940E",
        x"102F",
        x"5001",
        x"0911",
        x"3F08",
        x"EF8F",
        x"0718",
        x"F791",
        x"C002",
        x"940E",
        x"102F",
        x"9626",
        x"E0E4",
        x"940C",
        x"14F2",
        x"EF8F",
        x"BB87",
        x"E38F",
        x"BB81",
        x"B812",
        x"BA18",
        x"E020",
        x"EE31",
        x"E040",
        x"E050",
        x"E060",
        x"EE71",
        x"E080",
        x"E090",
        x"940E",
        x"146D",
        x"940E",
        x"0B5A",
        x"E060",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"047B",
        x"E060",
        x"E070",
        x"E08A",
        x"E090",
        x"940E",
        x"047B",
        x"E081",
        x"E090",
        x"940E",
        x"0D36",
        x"E061",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"0E2C",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E9EF",
        x"E1F1",
        x"940C",
        x"14D0",
        x"2EB8",
        x"2EA9",
        x"2F28",
        x"2F39",
        x"2F42",
        x"2F53",
        x"2EE4",
        x"2EF5",
        x"1AE2",
        x"0AF3",
        x"2F04",
        x"2F15",
        x"5F4F",
        x"4F5F",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"5681",
        x"318A",
        x"F390",
        x"EDE0",
        x"2ECE",
        x"E0E0",
        x"2EDE",
        x"E0C0",
        x"E0D0",
        x"2DEC",
        x"2DFD",
        x"9181",
        x"9191",
        x"2ECE",
        x"2EDF",
        x"2FE8",
        x"2FF9",
        x"9001",
        x"2000",
        x"F7E9",
        x"2F4E",
        x"2F5F",
        x"5041",
        x"0951",
        x"1B48",
        x"0B59",
        x"16E4",
        x"06F5",
        x"F414",
        x"2D4E",
        x"2D5F",
        x"2D6B",
        x"2D7A",
        x"940E",
        x"1569",
        x"2B89",
        x"F451",
        x"0FCC",
        x"1FDD",
        x"55CC",
        x"4FDF",
        x"81E8",
        x"81F9",
        x"2F80",
        x"2F91",
        x"9509",
        x"C016",
        x"9621",
        x"31C6",
        x"05D1",
        x"F6B1",
        x"92AF",
        x"92BF",
        x"E882",
        x"E090",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"14EC",
        x"E0A0",
        x"E0B0",
        x"E0E0",
        x"E1F2",
        x"940C",
        x"14C9",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"04AF",
        x"2F08",
        x"2F19",
        x"2FE8",
        x"2FF9",
        x"53EC",
        x"4FFB",
        x"95C8",
        x"2C30",
        x"2CE3",
        x"2CF1",
        x"E083",
        x"16E8",
        x"04F1",
        x"F06C",
        x"940E",
        x"04AF",
        x"2E78",
        x"2E69",
        x"E09C",
        x"16E9",
        x"04F1",
        x"F03C",
        x"940E",
        x"04AF",
        x"2E58",
        x"2E49",
        x"C004",
        x"2C71",
        x"2C61",
        x"2C51",
        x"2C41",
        x"2FE0",
        x"2FF1",
        x"53EC",
        x"4FFA",
        x"95C8",
        x"2D80",
        x"E090",
        x"E063",
        x"E070",
        x"940E",
        x"1490",
        x"2EE8",
        x"2EF9",
        x"93DF",
        x"93CF",
        x"EB8C",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E000",
        x"E010",
        x"2D8E",
        x"2D9F",
        x"538C",
        x"4F99",
        x"2EE8",
        x"2EF9",
        x"EB99",
        x"2E89",
        x"E094",
        x"2E99",
        x"E122",
        x"2EA2",
        x"E021",
        x"2EB2",
        x"2DEE",
        x"2DFF",
        x"0FE0",
        x"1FF1",
        x"95C8",
        x"2DE0",
        x"921F",
        x"93EF",
        x"929F",
        x"928F",
        x"E182",
        x"2EC8",
        x"E081",
        x"2ED8",
        x"92BF",
        x"92AF",
        x"940E",
        x"1579",
        x"5F0F",
        x"4F1F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"3003",
        x"0511",
        x"F719",
        x"EB87",
        x"E094",
        x"939F",
        x"938F",
        x"92DF",
        x"92CF",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2D43",
        x"E050",
        x"3141",
        x"0551",
        x"F008",
        x"C0CE",
        x"2FE4",
        x"2FF5",
        x"5DE0",
        x"4FFF",
        x"940C",
        x"1500",
        x"EA8E",
        x"E094",
        x"C002",
        x"EA85",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C0B6",
        x"2F2C",
        x"2F3D",
        x"5F2E",
        x"4F3F",
        x"0D27",
        x"1D31",
        x"FC77",
        x"953A",
        x"933F",
        x"932F",
        x"E98C",
        x"E094",
        x"C004",
        x"926F",
        x"927F",
        x"E981",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"9621",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"C095",
        x"926F",
        x"927F",
        x"E886",
        x"E094",
        x"CFEB",
        x"926F",
        x"927F",
        x"E78B",
        x"E094",
        x"CFE6",
        x"926F",
        x"927F",
        x"E780",
        x"E094",
        x"CFE1",
        x"926F",
        x"927F",
        x"E685",
        x"E094",
        x"CFDC",
        x"926F",
        x"927F",
        x"E58A",
        x"E094",
        x"CFD7",
        x"926F",
        x"927F",
        x"E48F",
        x"E094",
        x"CFD2",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"E482",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C05F",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"E385",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C047",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"E288",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C02F",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"E18B",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"C017",
        x"926F",
        x"927F",
        x"924F",
        x"925F",
        x"E08E",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"9622",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"E08C",
        x"E094",
        x"939F",
        x"938F",
        x"E182",
        x"E091",
        x"939F",
        x"938F",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"B7CD",
        x"B7DE",
        x"E1E1",
        x"940C",
        x"14E5",
        x"E0A0",
        x"E0B0",
        x"E6EB",
        x"E1F3",
        x"940C",
        x"14D0",
        x"E283",
        x"E090",
        x"940E",
        x"0494",
        x"2F08",
        x"2F19",
        x"E286",
        x"E090",
        x"940E",
        x"04BD",
        x"2EB8",
        x"2EA9",
        x"E284",
        x"E090",
        x"940E",
        x"04BD",
        x"2ED8",
        x"2EC9",
        x"E282",
        x"E090",
        x"940E",
        x"0494",
        x"2EF8",
        x"2EE9",
        x"E281",
        x"E090",
        x"940E",
        x"0494",
        x"2FC8",
        x"2FD9",
        x"E280",
        x"E090",
        x"940E",
        x"0494",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93DF",
        x"93CF",
        x"939F",
        x"938F",
        x"E98E",
        x"E097",
        x"939F",
        x"938F",
        x"E1C2",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"E983",
        x"E097",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"B78D",
        x"B79E",
        x"9642",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"EFCC",
        x"E0D0",
        x"E920",
        x"2EA2",
        x"E027",
        x"2EB2",
        x"E132",
        x"2EC3",
        x"E031",
        x"2ED3",
        x"FF07",
        x"C005",
        x"8188",
        x"2799",
        x"FD87",
        x"9590",
        x"C002",
        x"E28D",
        x"E090",
        x"939F",
        x"938F",
        x"92BF",
        x"92AF",
        x"E182",
        x"2EE8",
        x"E081",
        x"2EF8",
        x"92DF",
        x"92CF",
        x"940E",
        x"1579",
        x"0F00",
        x"1F11",
        x"9621",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"E091",
        x"30C4",
        x"07D9",
        x"F6F1",
        x"E88E",
        x"E097",
        x"939F",
        x"938F",
        x"92FF",
        x"92EF",
        x"940E",
        x"1579",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"14EC",
        x"93CF",
        x"93DF",
        x"EE89",
        x"E097",
        x"939F",
        x"938F",
        x"E0C4",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"EE82",
        x"E097",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"9508",
        x"93CF",
        x"93DF",
        x"3081",
        x"F419",
        x"940E",
        x"13EE",
        x"C01A",
        x"ED8D",
        x"E097",
        x"939F",
        x"938F",
        x"E1C2",
        x"E0D1",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"ED86",
        x"E097",
        x"939F",
        x"938F",
        x"93DF",
        x"93CF",
        x"940E",
        x"1579",
        x"B78D",
        x"B79E",
        x"9608",
        x"B60F",
        x"94F8",
        x"BF9E",
        x"BE0F",
        x"BF8D",
        x"91DF",
        x"91CF",
        x"9508",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"E188",
        x"B98A",
        x"EF67",
        x"E17E",
        x"E08F",
        x"E090",
        x"940E",
        x"14A1",
        x"5021",
        x"B929",
        x"9508",
        x"9508",
        x"9B5D",
        x"CFFE",
        x"B98C",
        x"9508",
        x"308D",
        x"F011",
        x"308A",
        x"F439",
        x"3061",
        x"F049",
        x"E08D",
        x"940E",
        x"1441",
        x"E08A",
        x"C002",
        x"3061",
        x"F011",
        x"940E",
        x"1441",
        x"9508",
        x"E060",
        x"940E",
        x"1445",
        x"E080",
        x"E090",
        x"9508",
        x"E061",
        x"940E",
        x"1445",
        x"E080",
        x"E090",
        x"9508",
        x"9508",
        x"9B5F",
        x"CFFE",
        x"B18C",
        x"9508",
        x"E080",
        x"9508",
        x"B18B",
        x"7880",
        x"9508",
        x"E080",
        x"9508",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F429",
        x"E188",
        x"B98A",
        x"E686",
        x"B989",
        x"C002",
        x"940E",
        x"1431",
        x"E080",
        x"940E",
        x"140D",
        x"940E",
        x"13EE",
        x"9508",
        x"9508",
        x"9508",
        x"940E",
        x"1170",
        x"E080",
        x"E090",
        x"940E",
        x"0D41",
        x"E180",
        x"E093",
        x"940E",
        x"0421",
        x"E180",
        x"E093",
        x"940E",
        x"1199",
        x"CFF7",
        x"2400",
        x"2755",
        x"C004",
        x"0E08",
        x"1F59",
        x"0F88",
        x"1F99",
        x"9700",
        x"F029",
        x"9576",
        x"9567",
        x"F3B8",
        x"0571",
        x"F7B9",
        x"2D80",
        x"2F95",
        x"9508",
        x"E2A1",
        x"2E1A",
        x"1BAA",
        x"1BBB",
        x"2FEA",
        x"2FFB",
        x"C00D",
        x"1FAA",
        x"1FBB",
        x"1FEE",
        x"1FFF",
        x"17A2",
        x"07B3",
        x"07E4",
        x"07F5",
        x"F020",
        x"1BA2",
        x"0BB3",
        x"0BE4",
        x"0BF5",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"941A",
        x"F769",
        x"9560",
        x"9570",
        x"9580",
        x"9590",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"1BCA",
        x"0BDB",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"9409",
        x"882A",
        x"8839",
        x"8848",
        x"845F",
        x"846E",
        x"847D",
        x"848C",
        x"849B",
        x"84AA",
        x"84B9",
        x"84C8",
        x"80DF",
        x"80EE",
        x"80FD",
        x"810C",
        x"811B",
        x"81AA",
        x"81B9",
        x"0FCE",
        x"1DD1",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2FCA",
        x"2FDB",
        x"9508",
        x"0FEE",
        x"1FFF",
        x"95C8",
        x"9631",
        x"920F",
        x"95C8",
        x"920F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E0EE",
        x"E1F5",
        x"940C",
        x"14CE",
        x"2FC8",
        x"2FD9",
        x"8168",
        x"8179",
        x"818A",
        x"819B",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F421",
        x"E264",
        x"ED79",
        x"E58B",
        x"E097",
        x"E12D",
        x"EF33",
        x"E041",
        x"E050",
        x"940E",
        x"1C0B",
        x"2E82",
        x"2E93",
        x"2EA4",
        x"2EB5",
        x"EA27",
        x"E431",
        x"E040",
        x"E050",
        x"940E",
        x"1C22",
        x"2EC2",
        x"2ED3",
        x"2EE4",
        x"2EF5",
        x"2D9B",
        x"2D8A",
        x"2D79",
        x"2D68",
        x"EE2C",
        x"EF34",
        x"EF4F",
        x"EF5F",
        x"940E",
        x"1C22",
        x"2F02",
        x"2F13",
        x"2F24",
        x"2F35",
        x"2DBF",
        x"2DAE",
        x"2D9D",
        x"2D8C",
        x"0F80",
        x"1F91",
        x"1FA2",
        x"1FB3",
        x"FFB7",
        x"C003",
        x"9701",
        x"09A1",
        x"48B0",
        x"8388",
        x"8399",
        x"83AA",
        x"83BB",
        x"779F",
        x"B7CD",
        x"B7DE",
        x"E0EC",
        x"940C",
        x"14EA",
        x"940E",
        x"1508",
        x"9508",
        x"E280",
        x"E091",
        x"940E",
        x"1508",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"9380",
        x"0120",
        x"9390",
        x"0121",
        x"93A0",
        x"0122",
        x"93B0",
        x"0123",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"5041",
        x"4050",
        x"F030",
        x"918D",
        x"9001",
        x"1980",
        x"F419",
        x"2000",
        x"F7B9",
        x"1B88",
        x"0B99",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E7EF",
        x"E1F5",
        x"940C",
        x"14D6",
        x"810F",
        x"8518",
        x"2FE0",
        x"2FF1",
        x"8183",
        x"6088",
        x"8383",
        x"2F4C",
        x"2F5D",
        x"5F45",
        x"4F5F",
        x"8569",
        x"857A",
        x"2F80",
        x"2F91",
        x"940E",
        x"15B3",
        x"2FE0",
        x"2FF1",
        x"8123",
        x"7F27",
        x"8323",
        x"E0E4",
        x"940C",
        x"14F2",
        x"E0AE",
        x"E0B0",
        x"E9EE",
        x"E1F5",
        x"940C",
        x"14D8",
        x"E085",
        x"838C",
        x"898B",
        x"899C",
        x"839A",
        x"8389",
        x"2F4C",
        x"2F5D",
        x"5E49",
        x"4F5F",
        x"896D",
        x"897E",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"196E",
        x"962E",
        x"E0E2",
        x"940C",
        x"14F4",
        x"E0AC",
        x"E0B0",
        x"EBE9",
        x"E1F5",
        x"940C",
        x"14C8",
        x"2EE8",
        x"2EF9",
        x"2EC6",
        x"2ED7",
        x"2F04",
        x"2F15",
        x"2FE8",
        x"2FF9",
        x"8217",
        x"8216",
        x"8183",
        x"FF81",
        x"C1EF",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2E88",
        x"2E99",
        x"2DEE",
        x"2DFF",
        x"8193",
        x"2DEC",
        x"2DFD",
        x"FD93",
        x"95C8",
        x"FF93",
        x"8000",
        x"9631",
        x"2D80",
        x"2ECE",
        x"2EDF",
        x"2388",
        x"F409",
        x"C1D5",
        x"3285",
        x"F451",
        x"FD93",
        x"95C8",
        x"FF93",
        x"8000",
        x"9631",
        x"2D80",
        x"2ECE",
        x"2EDF",
        x"3285",
        x"F431",
        x"2D6E",
        x"2D7F",
        x"E090",
        x"940E",
        x"1B4D",
        x"CFDE",
        x"2C51",
        x"2C31",
        x"E020",
        x"3220",
        x"F4A0",
        x"328B",
        x"F069",
        x"F430",
        x"3280",
        x"F059",
        x"3283",
        x"F469",
        x"6120",
        x"C02E",
        x"328D",
        x"F039",
        x"3380",
        x"F439",
        x"6021",
        x"C028",
        x"6022",
        x"6024",
        x"C025",
        x"6028",
        x"C023",
        x"FD27",
        x"C02E",
        x"ED30",
        x"0F38",
        x"303A",
        x"F488",
        x"FF26",
        x"C007",
        x"2D85",
        x"E06A",
        x"940E",
        x"1C02",
        x"2E58",
        x"0E53",
        x"C014",
        x"2D83",
        x"E06A",
        x"940E",
        x"1C02",
        x"2E38",
        x"0E33",
        x"6220",
        x"C00C",
        x"328E",
        x"F421",
        x"FD26",
        x"C18F",
        x"6420",
        x"C006",
        x"368C",
        x"F411",
        x"6820",
        x"C002",
        x"3688",
        x"F469",
        x"2DEC",
        x"2DFD",
        x"FD93",
        x"95C8",
        x"FF93",
        x"8000",
        x"9631",
        x"2D80",
        x"2ECE",
        x"2EDF",
        x"2388",
        x"F009",
        x"CFBA",
        x"2F98",
        x"7D9F",
        x"5495",
        x"3093",
        x"F428",
        x"5F0C",
        x"4F1F",
        x"E3FF",
        x"83F9",
        x"C00E",
        x"3683",
        x"F031",
        x"3783",
        x"F081",
        x"3583",
        x"F009",
        x"C06D",
        x"C029",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"8389",
        x"5F0E",
        x"4F1F",
        x"2444",
        x"9443",
        x"2C51",
        x"2CA8",
        x"2CB9",
        x"C01A",
        x"2E60",
        x"2E71",
        x"E0F2",
        x"0E6F",
        x"1C71",
        x"2FE0",
        x"2FF1",
        x"80A0",
        x"80B1",
        x"FF26",
        x"C003",
        x"2D65",
        x"E070",
        x"C002",
        x"EF6F",
        x"EF7F",
        x"2D8A",
        x"2D9B",
        x"872C",
        x"940E",
        x"1B02",
        x"2E48",
        x"2E59",
        x"2D06",
        x"2D17",
        x"852C",
        x"772F",
        x"2E22",
        x"C01C",
        x"2E60",
        x"2E71",
        x"E0F2",
        x"0E6F",
        x"1C71",
        x"2FE0",
        x"2FF1",
        x"80A0",
        x"80B1",
        x"FF26",
        x"C003",
        x"2D65",
        x"E070",
        x"C002",
        x"EF6F",
        x"EF7F",
        x"2D8A",
        x"2D9B",
        x"872C",
        x"940E",
        x"1AF5",
        x"2E48",
        x"2E59",
        x"852C",
        x"6820",
        x"2E22",
        x"2D06",
        x"2D17",
        x"FC23",
        x"C021",
        x"2D83",
        x"E090",
        x"1648",
        x"0659",
        x"F4E0",
        x"2D6E",
        x"2D7F",
        x"E280",
        x"E090",
        x"940E",
        x"1B4D",
        x"943A",
        x"CFF3",
        x"2DEA",
        x"2DFB",
        x"FC27",
        x"95C8",
        x"FE27",
        x"8000",
        x"9631",
        x"2D80",
        x"2EAE",
        x"2EBF",
        x"2D6E",
        x"2D7F",
        x"E090",
        x"940E",
        x"1B4D",
        x"1031",
        x"943A",
        x"E0F1",
        x"1A4F",
        x"0851",
        x"1441",
        x"0451",
        x"F749",
        x"C0F1",
        x"3684",
        x"F011",
        x"3689",
        x"F549",
        x"2FE0",
        x"2FF1",
        x"FF27",
        x"C007",
        x"8160",
        x"8171",
        x"8182",
        x"8193",
        x"5F0C",
        x"4F1F",
        x"C008",
        x"8160",
        x"8171",
        x"2788",
        x"FD77",
        x"9580",
        x"2F98",
        x"5F0E",
        x"4F1F",
        x"762F",
        x"2EB2",
        x"FF97",
        x"C009",
        x"9590",
        x"9580",
        x"9570",
        x"9561",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"6820",
        x"2EB2",
        x"E02A",
        x"E030",
        x"2D48",
        x"2D59",
        x"940E",
        x"1B9B",
        x"2EA8",
        x"18A8",
        x"C046",
        x"3785",
        x"F429",
        x"7E2F",
        x"2EB2",
        x"E02A",
        x"E030",
        x"C025",
        x"2FF2",
        x"7FF9",
        x"2EBF",
        x"368F",
        x"F0C1",
        x"F418",
        x"3588",
        x"F079",
        x"C0BF",
        x"3780",
        x"F019",
        x"3788",
        x"F021",
        x"C0BA",
        x"2F2F",
        x"6120",
        x"2EB2",
        x"FEB4",
        x"C00D",
        x"2D8B",
        x"6084",
        x"2EB8",
        x"C009",
        x"FF24",
        x"C00A",
        x"2F9F",
        x"6096",
        x"2EB9",
        x"C006",
        x"E028",
        x"E030",
        x"C005",
        x"E120",
        x"E030",
        x"C002",
        x"E120",
        x"E032",
        x"2FE0",
        x"2FF1",
        x"FEB7",
        x"C007",
        x"8160",
        x"8171",
        x"8182",
        x"8193",
        x"5F0C",
        x"4F1F",
        x"C006",
        x"8160",
        x"8171",
        x"E080",
        x"E090",
        x"5F0E",
        x"4F1F",
        x"2D48",
        x"2D59",
        x"940E",
        x"1B9B",
        x"2EA8",
        x"18A8",
        x"2DFB",
        x"77FF",
        x"2EBF",
        x"FEB6",
        x"C00B",
        x"2D2B",
        x"7F2E",
        x"14A5",
        x"F450",
        x"FEB4",
        x"C00A",
        x"FCB2",
        x"C008",
        x"2D2B",
        x"7E2E",
        x"C005",
        x"2C7A",
        x"2D2B",
        x"C003",
        x"2C7A",
        x"C001",
        x"2C75",
        x"FF24",
        x"C00E",
        x"2FEC",
        x"2FFD",
        x"0DEA",
        x"1DF1",
        x"8180",
        x"3380",
        x"F411",
        x"7E29",
        x"C009",
        x"FF22",
        x"C006",
        x"9473",
        x"9473",
        x"C004",
        x"2F82",
        x"7886",
        x"F009",
        x"9473",
        x"FD23",
        x"C014",
        x"FF20",
        x"C006",
        x"2C5A",
        x"1473",
        x"F418",
        x"0C53",
        x"1857",
        x"2C73",
        x"1473",
        x"F470",
        x"2D6E",
        x"2D7F",
        x"E280",
        x"E090",
        x"872C",
        x"940E",
        x"1B4D",
        x"9473",
        x"852C",
        x"CFF4",
        x"1473",
        x"F410",
        x"1837",
        x"C001",
        x"2C31",
        x"FF24",
        x"C014",
        x"2D6E",
        x"2D7F",
        x"E380",
        x"E090",
        x"872C",
        x"940E",
        x"1B4D",
        x"852C",
        x"FF22",
        x"C019",
        x"FF21",
        x"C003",
        x"E588",
        x"E090",
        x"C002",
        x"E788",
        x"E090",
        x"2D6E",
        x"2D7F",
        x"C00D",
        x"2F82",
        x"7886",
        x"F061",
        x"FD21",
        x"C002",
        x"E280",
        x"C001",
        x"E28B",
        x"FD27",
        x"E28D",
        x"2D6E",
        x"2D7F",
        x"E090",
        x"940E",
        x"1B4D",
        x"14A5",
        x"F440",
        x"2D6E",
        x"2D7F",
        x"E380",
        x"E090",
        x"940E",
        x"1B4D",
        x"945A",
        x"CFF6",
        x"94AA",
        x"2DE8",
        x"2DF9",
        x"0DEA",
        x"1DF1",
        x"8180",
        x"2D6E",
        x"2D7F",
        x"E090",
        x"940E",
        x"1B4D",
        x"20AA",
        x"F799",
        x"2033",
        x"F409",
        x"CE23",
        x"2D6E",
        x"2D7F",
        x"E280",
        x"E090",
        x"940E",
        x"1B4D",
        x"943A",
        x"CFF5",
        x"2DEE",
        x"2DFF",
        x"8186",
        x"8197",
        x"C002",
        x"EF8F",
        x"EF9F",
        x"962C",
        x"E1E2",
        x"940C",
        x"14E4",
        x"FD20",
        x"C00A",
        x"2FE8",
        x"2FF9",
        x"FD23",
        x"C005",
        x"FF22",
        x"C002",
        x"8373",
        x"8362",
        x"8351",
        x"8340",
        x"9508",
        x"FD44",
        x"C012",
        x"FD46",
        x"C012",
        x"2FA6",
        x"2FB7",
        x"2FE8",
        x"2FF9",
        x"0FAA",
        x"1FBB",
        x"1FEE",
        x"1FFF",
        x"9410",
        x"F7D1",
        x"0F6A",
        x"1F7B",
        x"1F8E",
        x"1F9F",
        x"E031",
        x"C003",
        x"E033",
        x"C001",
        x"E034",
        x"0F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"5031",
        x"F7D1",
        x"0F62",
        x"1D71",
        x"1D81",
        x"1D91",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"2F80",
        x"2F91",
        x"940E",
        x"1B0E",
        x"2FC8",
        x"2FD9",
        x"FD97",
        x"C00A",
        x"940E",
        x"1ADE",
        x"2B89",
        x"F7A1",
        x"2F60",
        x"2F71",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1B81",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2EA6",
        x"2E84",
        x"2E95",
        x"2F02",
        x"940E",
        x"1B0E",
        x"2F48",
        x"2F59",
        x"2755",
        x"324B",
        x"0551",
        x"F021",
        x"324D",
        x"0551",
        x"F459",
        x"6800",
        x"94AA",
        x"F411",
        x"E080",
        x"C075",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1B0E",
        x"FD97",
        x"CFF8",
        x"2F10",
        x"7F1D",
        x"2F30",
        x"7330",
        x"F511",
        x"3380",
        x"F501",
        x"24FF",
        x"94FA",
        x"0CFA",
        x"F409",
        x"C04B",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1B0E",
        x"FD97",
        x"C045",
        x"2F38",
        x"7D3F",
        x"3538",
        x"F459",
        x"6412",
        x"94AA",
        x"94AA",
        x"F1E9",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1B0E",
        x"FF97",
        x"C007",
        x"C036",
        x"FF06",
        x"C002",
        x"6012",
        x"C001",
        x"6112",
        x"2CAF",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"ED20",
        x"0F28",
        x"3028",
        x"F088",
        x"FF14",
        x"C005",
        x"2F6C",
        x"2F7D",
        x"940E",
        x"1B81",
        x"C01E",
        x"302A",
        x"F040",
        x"FF16",
        x"CFF7",
        x"7D2F",
        x"EE3F",
        x"0F32",
        x"3036",
        x"F790",
        x"5027",
        x"2F41",
        x"2D9F",
        x"2D8E",
        x"2D7D",
        x"2D6C",
        x"940E",
        x"17C8",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"6012",
        x"94AA",
        x"F069",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1B0E",
        x"FF97",
        x"CFD7",
        x"FD11",
        x"C005",
        x"CFA1",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"FF17",
        x"C008",
        x"94F0",
        x"94E0",
        x"94D0",
        x"94C0",
        x"1CC1",
        x"1CD1",
        x"1CE1",
        x"1CF1",
        x"2F21",
        x"2D7F",
        x"2D6E",
        x"2D5D",
        x"2D4C",
        x"2D88",
        x"2D99",
        x"940E",
        x"17BB",
        x"E081",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"E2A1",
        x"E0B0",
        x"EBE1",
        x"E1F8",
        x"940C",
        x"14CD",
        x"2EA8",
        x"2EB9",
        x"2EE4",
        x"2EF5",
        x"2F0C",
        x"2F1D",
        x"5F0F",
        x"4F1F",
        x"2EC0",
        x"2ED1",
        x"E280",
        x"2FA0",
        x"2FB1",
        x"921D",
        x"958A",
        x"F7E9",
        x"2DEA",
        x"2DFB",
        x"8073",
        x"E040",
        x"E050",
        x"2C81",
        x"E0B0",
        x"2C91",
        x"E081",
        x"E090",
        x"2FE2",
        x"2FF3",
        x"FC73",
        x"95C8",
        x"FE73",
        x"8000",
        x"9631",
        x"2DA0",
        x"2F0E",
        x"2F1F",
        x"2F7A",
        x"2F2E",
        x"2F3F",
        x"23AA",
        x"F419",
        x"E080",
        x"E090",
        x"C08D",
        x"35AE",
        x"F419",
        x"1541",
        x"0551",
        x"F179",
        x"2DE9",
        x"E0F0",
        x"17E4",
        x"07F5",
        x"F43C",
        x"35AD",
        x"F189",
        x"32AD",
        x"F419",
        x"23BB",
        x"F139",
        x"C003",
        x"23BB",
        x"F409",
        x"2E8A",
        x"2FE7",
        x"95E6",
        x"95E6",
        x"95E6",
        x"2D0C",
        x"2D1D",
        x"0F0E",
        x"1D11",
        x"2FE0",
        x"2FF1",
        x"2FA7",
        x"70A7",
        x"2F08",
        x"2F19",
        x"C002",
        x"0F00",
        x"1F11",
        x"95AA",
        x"F7E2",
        x"2FA0",
        x"2FB1",
        x"81B0",
        x"2BBA",
        x"83B0",
        x"1578",
        x"F059",
        x"1578",
        x"F410",
        x"5F7F",
        x"CFE2",
        x"5071",
        x"CFE0",
        x"2499",
        x"9493",
        x"C003",
        x"E0B1",
        x"C001",
        x"E0B0",
        x"5F4F",
        x"4F5F",
        x"CFB1",
        x"23BB",
        x"F019",
        x"818E",
        x"6280",
        x"838E",
        x"2099",
        x"F419",
        x"2499",
        x"9493",
        x"C01A",
        x"2DEC",
        x"2DFD",
        x"2F8C",
        x"2F9D",
        x"9681",
        x"8120",
        x"9520",
        x"9321",
        x"17E8",
        x"07F9",
        x"F7D1",
        x"CFF1",
        x"14E1",
        x"04F1",
        x"F041",
        x"2DAE",
        x"2DBF",
        x"938C",
        x"2DEE",
        x"2DFF",
        x"9631",
        x"2EEE",
        x"2EFF",
        x"5061",
        x"F129",
        x"2C91",
        x"2D8A",
        x"2D9B",
        x"A369",
        x"940E",
        x"1B0E",
        x"A169",
        x"FD97",
        x"C019",
        x"2F28",
        x"9526",
        x"9526",
        x"9526",
        x"2DEC",
        x"2DFD",
        x"0FE2",
        x"1DF1",
        x"8120",
        x"E030",
        x"2F48",
        x"2F59",
        x"7047",
        x"2755",
        x"C002",
        x"9535",
        x"9527",
        x"954A",
        x"F7E2",
        x"FD20",
        x"CFD5",
        x"2D6A",
        x"2D7B",
        x"940E",
        x"1B81",
        x"2099",
        x"F009",
        x"CF78",
        x"14E1",
        x"04F1",
        x"F019",
        x"2DAE",
        x"2DBF",
        x"921C",
        x"2F80",
        x"2F91",
        x"96A1",
        x"E0ED",
        x"940C",
        x"14E9",
        x"924F",
        x"925F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"921F",
        x"B7CD",
        x"B7DE",
        x"2F08",
        x"2F19",
        x"2E46",
        x"2E57",
        x"2EE4",
        x"2EF5",
        x"2FE8",
        x"2FF9",
        x"8217",
        x"8216",
        x"2CA1",
        x"2FE0",
        x"2FF1",
        x"80D3",
        x"2DE4",
        x"2DF5",
        x"FCD3",
        x"95C8",
        x"FED3",
        x"8000",
        x"9631",
        x"2D80",
        x"2F38",
        x"2E4E",
        x"2E5F",
        x"2388",
        x"F409",
        x"C12C",
        x"E090",
        x"8339",
        x"940E",
        x"1ADE",
        x"8139",
        x"2B89",
        x"F029",
        x"2F80",
        x"2F91",
        x"940E",
        x"17EA",
        x"CFE3",
        x"3235",
        x"F461",
        x"2DE4",
        x"2DF5",
        x"FCD3",
        x"95C8",
        x"FED3",
        x"8000",
        x"9631",
        x"2D30",
        x"2E4E",
        x"2E5F",
        x"3235",
        x"F481",
        x"2F80",
        x"2F91",
        x"8339",
        x"940E",
        x"1B0E",
        x"8139",
        x"FD97",
        x"C108",
        x"1738",
        x"F409",
        x"CFCA",
        x"2F60",
        x"2F71",
        x"940E",
        x"1B81",
        x"C102",
        x"323A",
        x"F459",
        x"FCD3",
        x"95C8",
        x"FED3",
        x"8000",
        x"9631",
        x"2D30",
        x"2E4E",
        x"2E5F",
        x"24BB",
        x"94B3",
        x"C001",
        x"2CB1",
        x"2C71",
        x"ED20",
        x"0F23",
        x"302A",
        x"F4B0",
        x"2DFB",
        x"60F2",
        x"2EBF",
        x"2D67",
        x"E070",
        x"E080",
        x"E090",
        x"E240",
        x"940E",
        x"17C8",
        x"2E76",
        x"2DE4",
        x"2DF5",
        x"FCD3",
        x"95C8",
        x"FED3",
        x"8000",
        x"9631",
        x"2D30",
        x"2E4E",
        x"2E5F",
        x"CFE6",
        x"FEB1",
        x"C003",
        x"2077",
        x"F419",
        x"C0D4",
        x"2477",
        x"947A",
        x"3638",
        x"F019",
        x"363C",
        x"F081",
        x"C01C",
        x"2DE4",
        x"2DF5",
        x"FCD3",
        x"95C8",
        x"FED3",
        x"8000",
        x"9631",
        x"2D30",
        x"2E4E",
        x"2E5F",
        x"3638",
        x"F481",
        x"2DFB",
        x"60F8",
        x"2EBF",
        x"2D8B",
        x"6084",
        x"2EB8",
        x"2DE4",
        x"2DF5",
        x"FCD3",
        x"95C8",
        x"FED3",
        x"8000",
        x"9631",
        x"2D30",
        x"2E4E",
        x"2E5F",
        x"2333",
        x"F409",
        x"C0AE",
        x"2F63",
        x"E070",
        x"EE8E",
        x"E097",
        x"8339",
        x"940E",
        x"1AE6",
        x"8139",
        x"2B89",
        x"F409",
        x"C0A3",
        x"FCB0",
        x"C00A",
        x"2DEE",
        x"2DFF",
        x"80C0",
        x"80D1",
        x"2D8E",
        x"2D9F",
        x"9602",
        x"2EE8",
        x"2EF9",
        x"C002",
        x"2CC1",
        x"2CD1",
        x"363E",
        x"F461",
        x"2FE0",
        x"2FF1",
        x"8146",
        x"8157",
        x"E060",
        x"E070",
        x"2D2B",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"17BB",
        x"CF4A",
        x"3633",
        x"F4C1",
        x"FCB1",
        x"C002",
        x"2477",
        x"9473",
        x"2F80",
        x"2F91",
        x"940E",
        x"1B0E",
        x"FD97",
        x"C079",
        x"14C1",
        x"04D1",
        x"F041",
        x"2DEC",
        x"2DFD",
        x"8380",
        x"2D8C",
        x"2D9D",
        x"9601",
        x"2EC8",
        x"2ED9",
        x"947A",
        x"F769",
        x"C067",
        x"353B",
        x"F479",
        x"2D24",
        x"2D35",
        x"2D4C",
        x"2D5D",
        x"2D67",
        x"2F80",
        x"2F91",
        x"940E",
        x"18AB",
        x"2E48",
        x"2E59",
        x"9700",
        x"F009",
        x"C057",
        x"C050",
        x"2F80",
        x"2F91",
        x"8339",
        x"940E",
        x"17EA",
        x"8139",
        x"FD97",
        x"C052",
        x"363F",
        x"F1A9",
        x"F428",
        x"3634",
        x"F171",
        x"3639",
        x"F1B9",
        x"C033",
        x"3733",
        x"F081",
        x"3735",
        x"F139",
        x"C02E",
        x"14C1",
        x"04D1",
        x"F041",
        x"2DEC",
        x"2DFD",
        x"8280",
        x"2D8C",
        x"2D9D",
        x"9601",
        x"2EC8",
        x"2ED9",
        x"947A",
        x"F091",
        x"2F80",
        x"2F91",
        x"940E",
        x"1B0E",
        x"2E88",
        x"2E99",
        x"FD97",
        x"C00A",
        x"940E",
        x"1ADE",
        x"2B89",
        x"F339",
        x"2F60",
        x"2F71",
        x"2D88",
        x"2D99",
        x"940E",
        x"1B81",
        x"14C1",
        x"04D1",
        x"F0F9",
        x"2DEC",
        x"2DFD",
        x"8210",
        x"C01B",
        x"2DFB",
        x"62F0",
        x"2EBF",
        x"C007",
        x"2D8B",
        x"6180",
        x"2EB8",
        x"C003",
        x"2D9B",
        x"6490",
        x"2EB9",
        x"2D2B",
        x"2D4C",
        x"2D5D",
        x"2D67",
        x"2F80",
        x"2F91",
        x"940E",
        x"1809",
        x"2388",
        x"F431",
        x"2FE0",
        x"2FF1",
        x"8183",
        x"7380",
        x"F429",
        x"C006",
        x"FCB0",
        x"CEC7",
        x"94A3",
        x"CEC5",
        x"20AA",
        x"F019",
        x"2D8A",
        x"E090",
        x"C002",
        x"EF8F",
        x"EF9F",
        x"900F",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"907F",
        x"905F",
        x"904F",
        x"9508",
        x"1191",
        x"C11F",
        x"3280",
        x"F019",
        x"5089",
        x"5085",
        x"F7D0",
        x"9508",
        x"2FE8",
        x"2FF9",
        x"95C8",
        x"9631",
        x"1606",
        x"F029",
        x"2000",
        x"F7D1",
        x"2D80",
        x"2D91",
        x"9508",
        x"9731",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"2FE8",
        x"2FF9",
        x"95C8",
        x"9631",
        x"5061",
        x"4070",
        x"1001",
        x"F7D0",
        x"9580",
        x"9590",
        x"0F8E",
        x"1F9F",
        x"9508",
        x"2FE8",
        x"2FF9",
        x"5061",
        x"4070",
        x"9001",
        x"1001",
        x"F7D8",
        x"9580",
        x"9590",
        x"0F8E",
        x"1F9F",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"812B",
        x"FF20",
        x"C033",
        x"FF26",
        x"C00A",
        x"7B2F",
        x"832B",
        x"818E",
        x"819F",
        x"9601",
        x"839F",
        x"838E",
        x"818A",
        x"E090",
        x"C029",
        x"FF22",
        x"C00F",
        x"81E8",
        x"81F9",
        x"8180",
        x"2799",
        x"FD87",
        x"9590",
        x"9700",
        x"F419",
        x"6220",
        x"832B",
        x"C01A",
        x"9631",
        x"83F9",
        x"83E8",
        x"C00E",
        x"85EA",
        x"85FB",
        x"9509",
        x"FF97",
        x"C009",
        x"812B",
        x"9601",
        x"F411",
        x"E180",
        x"C001",
        x"E280",
        x"2B82",
        x"838B",
        x"C008",
        x"812E",
        x"813F",
        x"5F2F",
        x"4F3F",
        x"833F",
        x"832E",
        x"2799",
        x"C002",
        x"EF8F",
        x"EF9F",
        x"91DF",
        x"91CF",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F18",
        x"2F09",
        x"2FC6",
        x"2FD7",
        x"818B",
        x"FD81",
        x"C003",
        x"EF8F",
        x"EF9F",
        x"C021",
        x"FF82",
        x"C011",
        x"814E",
        x"815F",
        x"812C",
        x"813D",
        x"1742",
        x"0753",
        x"F484",
        x"81E8",
        x"81F9",
        x"2F2E",
        x"2F3F",
        x"5F2F",
        x"4F3F",
        x"8339",
        x"8328",
        x"8310",
        x"C006",
        x"85E8",
        x"85F9",
        x"2F81",
        x"9509",
        x"2B89",
        x"F721",
        x"812E",
        x"813F",
        x"5F2F",
        x"4F3F",
        x"833F",
        x"832E",
        x"2F81",
        x"2F90",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"8123",
        x"FF20",
        x"C012",
        x"FD26",
        x"C010",
        x"3F8F",
        x"EF3F",
        x"0793",
        x"F061",
        x"8382",
        x"7D2F",
        x"6420",
        x"8323",
        x"8126",
        x"8137",
        x"5021",
        x"0931",
        x"8337",
        x"8326",
        x"2799",
        x"9508",
        x"EF8F",
        x"EF9F",
        x"9508",
        x"2FE4",
        x"2FF5",
        x"27AA",
        x"3028",
        x"F169",
        x"3120",
        x"F199",
        x"94E8",
        x"936F",
        x"7F6E",
        x"5F6E",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"4FAF",
        x"E0B1",
        x"D041",
        x"E0B4",
        x"D03F",
        x"0F67",
        x"1F78",
        x"1F89",
        x"1F9A",
        x"1DA1",
        x"0F68",
        x"1F79",
        x"1F8A",
        x"1D91",
        x"1DA1",
        x"0F6A",
        x"1D71",
        x"1D81",
        x"1D91",
        x"1DA1",
        x"D023",
        x"F409",
        x"9468",
        x"913F",
        x"2E06",
        x"0C00",
        x"1930",
        x"0C00",
        x"0C00",
        x"1930",
        x"5D30",
        x"9331",
        x"F6CE",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"2F46",
        x"7047",
        x"5D40",
        x"9341",
        x"E0B3",
        x"D00F",
        x"F7C9",
        x"CFF5",
        x"2F46",
        x"704F",
        x"5D40",
        x"334A",
        x"F018",
        x"5D49",
        x"FD31",
        x"5240",
        x"9341",
        x"D002",
        x"F7A9",
        x"CFE9",
        x"E0B4",
        x"95A6",
        x"9597",
        x"9587",
        x"9577",
        x"9567",
        x"95BA",
        x"F7C9",
        x"9700",
        x"0561",
        x"0571",
        x"9508",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"2E0A",
        x"9406",
        x"9557",
        x"9547",
        x"9537",
        x"9527",
        x"95BA",
        x"F7C9",
        x"0F62",
        x"1F73",
        x"1F84",
        x"1F95",
        x"1DA0",
        x"9508",
        x"2799",
        x"2788",
        x"9508",
        x"2400",
        x"FD80",
        x"0E06",
        x"0F66",
        x"F011",
        x"9586",
        x"F7D1",
        x"2D80",
        x"9508",
        x"2E05",
        x"FB97",
        x"F41E",
        x"9400",
        x"940E",
        x"1C48",
        x"FD57",
        x"D007",
        x"940E",
        x"14A1",
        x"FC07",
        x"D003",
        x"F44E",
        x"940C",
        x"1C48",
        x"9550",
        x"9540",
        x"9530",
        x"9521",
        x"4F3F",
        x"4F4F",
        x"4F5F",
        x"9508",
        x"9468",
        x"1000",
        x"94E8",
        x"E0A0",
        x"E0B0",
        x"E2EB",
        x"E1FC",
        x"940C",
        x"14D0",
        x"EFEF",
        x"F9E7",
        x"2EA2",
        x"2EB3",
        x"2EC4",
        x"2ED5",
        x"235E",
        x"0F55",
        x"08EE",
        x"2CFE",
        x"2D0E",
        x"2D1F",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"239E",
        x"0F99",
        x"0B66",
        x"2F76",
        x"2F86",
        x"2F97",
        x"940E",
        x"1C50",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"14EC",
        x"9590",
        x"9580",
        x"9570",
        x"9561",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"9508",
        x"93DF",
        x"93CF",
        x"929F",
        x"E4A0",
        x"2E9A",
        x"2400",
        x"2DA0",
        x"2DB1",
        x"2DC0",
        x"2DD1",
        x"2DE0",
        x"2DF1",
        x"9516",
        x"9507",
        x"94F7",
        x"94E7",
        x"94D7",
        x"94C7",
        x"94B7",
        x"94A7",
        x"F448",
        x"6810",
        x"0FA2",
        x"1FB3",
        x"1FC4",
        x"1FD5",
        x"1FE6",
        x"1FF7",
        x"1E08",
        x"1E19",
        x"0F22",
        x"1F33",
        x"1F44",
        x"1F55",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"949A",
        x"F721",
        x"2F2A",
        x"2F3B",
        x"2F4C",
        x"2F5D",
        x"2F6E",
        x"2F7F",
        x"2D80",
        x"2D91",
        x"2411",
        x"909F",
        x"91CF",
        x"91DF",
        x"9508",
        x"94F8",
        x"CFFF",
        x"0001",
        x"0000",
        x"0169",
        x"016F",
        x"017C",
        x"0191",
        x"01A1",
        x"01B9",
        x"01C0",
        x"01C6",
        x"01C7",
        x"01CE",
        x"01D2",
        x"01DD",
        x"01E1",
        x"01EB",
        x"01D3",
        x"01F6",
        x"01DE",
        x"01EC",
        x"01DA",
        x"0201",
        x"0202",
        x"020B",
        x"0212",
        x"021F",
        x"022C",
        x"0239",
        x"0246",
        x"0252",
        x"025E",
        x"026A",
        x"0276",
        x"027F",
        x"0B94",
        x"0D41",
        x"1365",
        x"0548",
        x"0617",
        x"0574",
        x"0798",
        x"0884",
        x"0803",
        x"1112",
        x"0B22",
        x"0A77",
        x"0E5F",
        x"093B",
        x"0FDF",
        x"0FE4",
        x"0FE9",
        x"0FEE",
        x"0FF3",
        x"0FF8",
        x"0C21",
        x"0CB7",
        x"0288",
        x"028D",
        x"0296",
        x"029B",
        x"029F",
        x"02A4",
        x"02A8",
        x"02AC",
        x"02B0",
        x"02B4",
        x"02B9",
        x"02BF",
        x"02C4",
        x"02CA",
        x"02D0",
        x"02D7",
        x"02DE",
        x"02E6",
        x"02EE",
        x"02F6",
        x"02FE",
        x"0304",
        x"564E",
        x"422D",
        x"4944",
        x"435A",
        x"0000",
        x"0200",
        x"0000",
        x"0000",
        x"145B",
        x"0000",
        x"0000",
        x"0000",
        x"0200",
        x"0000",
        x"0000",
        x"1455",
        x"0000",
        x"0000",
        x"0001",
        x"0000",
        x"7825",
        x"2520",
        x"2078",
        x"7825",
        x"2500",
        x"2078",
        x"7825",
        x"2520",
        x"646C",
        x"3000",
        x"372E",
        x"0032",
        x"4349",
        x"2D45",
        x"3654",
        x"0035",
        x"6F4E",
        x"2076",
        x"3631",
        x"3220",
        x"3130",
        x"0035",
        x"3232",
        x"303A",
        x"3A33",
        x"3231",
        x"2500",
        x"782A",
        x"2520",
        x"0078",
        x"7825",
        x"2520",
        x"2078",
        x"6425",
        x"4600",
        x"7869",
        x"6465",
        x"4300",
        x"6568",
        x"6B63",
        x"7265",
        x"6F62",
        x"7261",
        x"0064",
        x"6E49",
        x"6576",
        x"7372",
        x"2065",
        x"6863",
        x"6365",
        x"656B",
        x"6272",
        x"616F",
        x"6472",
        x"4100",
        x"6464",
        x"6572",
        x"7373",
        x"7020",
        x"7461",
        x"6574",
        x"6E72",
        x"4900",
        x"766E",
        x"7265",
        x"6573",
        x"6120",
        x"6464",
        x"6572",
        x"7373",
        x"7020",
        x"7461",
        x"6574",
        x"6E72",
        x"5200",
        x"6E61",
        x"6F64",
        x"006D",
        x"654E",
        x"6576",
        x"0072",
        x"547E",
        x"2030",
        x"6E61",
        x"2064",
        x"547E",
        x"0031",
        x"547E",
        x"2030",
        x"6E61",
        x"2064",
        x"3154",
        x"7E00",
        x"3054",
        x"5400",
        x"2030",
        x"6F78",
        x"2072",
        x"3154",
        x"7E00",
        x"3054",
        x"6F20",
        x"2072",
        x"547E",
        x"0031",
        x"3054",
        x"7820",
        x"6F6E",
        x"2072",
        x"3154",
        x"7E00",
        x"3054",
        x"6F20",
        x"2072",
        x"3154",
        x"4100",
        x"776C",
        x"7961",
        x"0073",
        x"654D",
        x"206D",
        x"6452",
        x"4220",
        x"6B72",
        x"7470",
        x"4D00",
        x"6D65",
        x"5220",
        x"2064",
        x"6157",
        x"6374",
        x"0068",
        x"654D",
        x"206D",
        x"7257",
        x"4220",
        x"6B72",
        x"7470",
        x"4D00",
        x"6D65",
        x"5720",
        x"2072",
        x"6157",
        x"6374",
        x"0068",
        x"4F49",
        x"5220",
        x"2064",
        x"7242",
        x"706B",
        x"0074",
        x"4F49",
        x"5220",
        x"2064",
        x"6157",
        x"6374",
        x"0068",
        x"4F49",
        x"5720",
        x"2072",
        x"7242",
        x"706B",
        x"0074",
        x"4F49",
        x"5720",
        x"2072",
        x"6157",
        x"6374",
        x"0068",
        x"7845",
        x"4220",
        x"6B72",
        x"7470",
        x"4500",
        x"2078",
        x"6157",
        x"6374",
        x"0068",
        x"6568",
        x"706C",
        x"6300",
        x"6E6F",
        x"6974",
        x"756E",
        x"0065",
        x"6572",
        x"7367",
        x"6400",
        x"7369",
        x"6600",
        x"6C69",
        x"006C",
        x"7263",
        x"0063",
        x"656D",
        x"006D",
        x"6472",
        x"006D",
        x"7277",
        x"006D",
        x"6574",
        x"7473",
        x"7200",
        x"7365",
        x"7465",
        x"7300",
        x"6574",
        x"0070",
        x"7274",
        x"6361",
        x"0065",
        x"6C62",
        x"7369",
        x"0074",
        x"7262",
        x"6165",
        x"786B",
        x"7700",
        x"7461",
        x"6863",
        x"0078",
        x"7262",
        x"6165",
        x"726B",
        x"006D",
        x"6177",
        x"6374",
        x"7268",
        x"006D",
        x"7262",
        x"6165",
        x"776B",
        x"006D",
        x"6177",
        x"6374",
        x"7768",
        x"006D",
        x"6C63",
        x"6165",
        x"0072",
        x"7274",
        x"6769",
        x"6567",
        x"0072",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000"
    );

begin

    process (cp2)
    begin
        if rising_edge(cp2) then
            if ce = '1' then
                if (we = '1') then
                    RAM(conv_integer(address)) <= din;
                end if;
                dout <= RAM(conv_integer(address));
            end if;
        end if;
    end process;

end RTL;

