library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

-- This contains 0.986 of the ICE-65C02 firmware

-- For f_log2 definition
use WORK.SynthCtrlPack.all;

entity XPM is
    generic (
        WIDTH : integer;
        SIZE  : integer
    );
    port(
        cp2     : in  std_logic;
        ce      : in  std_logic;
        address : in  std_logic_vector(f_log2(SIZE) - 1 downto 0);
        din     : in  std_logic_vector(WIDTH - 1 downto 0);
        dout    : out std_logic_vector(WIDTH - 1 downto 0);
        we      : in  std_logic
    );
end;

architecture RTL of XPM is

    type ram_type is array (0 to SIZE - 1) of std_logic_vector (WIDTH - 1 downto 0);

    signal RAM : ram_type := (
        x"940C",
        x"0557",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"940C",
        x"0579",
        x"18A4",
        x"1970",
        x"18AA",
        x"18B8",
        x"18BE",
        x"18CC",
        x"18DD",
        x"18ED",
        x"18F6",
        x"18E4",
        x"1970",
        x"190D",
        x"1917",
        x"1929",
        x"193F",
        x"1954",
        x"205D",
        x"2000",
        x"2A2A",
        x"0A2A",
        x"6D00",
        x"6D65",
        x"726F",
        x"2079",
        x"6974",
        x"656D",
        x"756F",
        x"0074",
        x"696D",
        x"7373",
        x"6E69",
        x"2067",
        x"6C63",
        x"636F",
        x"006B",
        x"2A2A",
        x"202A",
        x"4900",
        x"746E",
        x"7265",
        x"7572",
        x"7470",
        x"6465",
        x"000A",
        x"5043",
        x"2055",
        x"7266",
        x"6565",
        x"7220",
        x"6E75",
        x"696E",
        x"676E",
        x"2E2E",
        x"0A2E",
        x"2000",
        x"203D",
        x"2000",
        x"2020",
        x"0020",
        x"7254",
        x"6769",
        x"6567",
        x"2072",
        x"6F43",
        x"6564",
        x"3A73",
        x"000A",
        x"6120",
        x"2074",
        x"5200",
        x"6D65",
        x"766F",
        x"6E69",
        x"2067",
        x"4E00",
        x"206F",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"6573",
        x"0A74",
        x"2900",
        x"000A",
        x"203A",
        x"2000",
        x"616D",
        x"6B73",
        x"0020",
        x"203A",
        x"2000",
        x"6E65",
        x"6261",
        x"656C",
        x"0A64",
        x"2000",
        x"6E69",
        x"6968",
        x"6962",
        x"6574",
        x"0A64",
        x"7300",
        x"696B",
        x"7070",
        x"6E69",
        x"2067",
        x"0053",
        x"2D20",
        x"3020",
        x"0078",
        x"6220",
        x"7479",
        x"7365",
        x"7420",
        x"206F",
        x"7830",
        x"7400",
        x"6172",
        x"736E",
        x"6566",
        x"7272",
        x"6465",
        x"3020",
        x"0078",
        x"6220",
        x"6461",
        x"7220",
        x"6365",
        x"726F",
        x"7364",
        x"000A",
        x"6720",
        x"6F6F",
        x"2064",
        x"6572",
        x"6F63",
        x"6472",
        x"2C73",
        x"0020",
        x"6572",
        x"6563",
        x"7669",
        x"6465",
        x"0020",
        x"7420",
        x"206F",
        x"5700",
        x"6F72",
        x"6574",
        x"0020",
        x"7250",
        x"7365",
        x"2073",
        x"6E61",
        x"2079",
        x"656B",
        x"2079",
        x"6F74",
        x"7320",
        x"6174",
        x"7472",
        x"7420",
        x"6172",
        x"736E",
        x"696D",
        x"7373",
        x"6F69",
        x"206E",
        x"6128",
        x"646E",
        x"6120",
        x"6167",
        x"6E69",
        x"6120",
        x"2074",
        x"6E65",
        x"2964",
        x"000A",
        x"2F20",
        x"003D",
        x"6F43",
        x"706D",
        x"7261",
        x"2065",
        x"6166",
        x"6C69",
        x"6465",
        x"003A",
        x"7263",
        x"3A63",
        x"0020",
        x"3D20",
        x"0020",
        x"7420",
        x"206F",
        x"5700",
        x"3A72",
        x"0020",
        x"6C46",
        x"7375",
        x"6968",
        x"676E",
        x"4520",
        x"6576",
        x"746E",
        x"4620",
        x"4649",
        x"0A4F",
        x"2000",
        x"6E69",
        x"7473",
        x"7572",
        x"7463",
        x"6F69",
        x"736E",
        x"000A",
        x"6E49",
        x"6574",
        x"7272",
        x"7075",
        x"6574",
        x"2064",
        x"6661",
        x"6574",
        x"2072",
        x"2000",
        x"6E69",
        x"7473",
        x"7572",
        x"7463",
        x"6F69",
        x"736E",
        x"000A",
        x"7453",
        x"7065",
        x"6970",
        x"676E",
        x"0020",
        x"754E",
        x"626D",
        x"7265",
        x"6F20",
        x"2066",
        x"6E69",
        x"7473",
        x"6375",
        x"6974",
        x"6E6F",
        x"2073",
        x"756D",
        x"7473",
        x"6220",
        x"2065",
        x"6F70",
        x"6973",
        x"6974",
        x"6576",
        x"000A",
        x"6F43",
        x"6D6D",
        x"6E61",
        x"7364",
        x"0A3A",
        x"2000",
        x"2020",
        x"5200",
        x"7365",
        x"7465",
        x"6974",
        x"676E",
        x"4320",
        x"5550",
        x"000A",
        x"203A",
        x"6170",
        x"7373",
        x"6465",
        x"000A",
        x"6520",
        x"7272",
        x"726F",
        x"0A73",
        x"3A00",
        x"6620",
        x"6961",
        x"656C",
        x"3A64",
        x"0020",
        x"654D",
        x"6F6D",
        x"7972",
        x"7420",
        x"7365",
        x"3A74",
        x"0020",
        x"0A29",
        x"2C00",
        x"5220",
        x"6165",
        x"2064",
        x"6162",
        x"6B63",
        x"0020",
        x"2820",
        x"7257",
        x"746F",
        x"3A65",
        x"0020",
        x"6146",
        x"6C69",
        x"6120",
        x"2074",
        x"2000",
        x"6C61",
        x"6572",
        x"6461",
        x"2079",
        x"6573",
        x"2074",
        x"7461",
        x"0020",
        x"6220",
        x"6572",
        x"6B61",
        x"6F70",
        x"6E69",
        x"7374",
        x"6120",
        x"6572",
        x"6120",
        x"726C",
        x"6165",
        x"7964",
        x"7320",
        x"7465",
        x"000A",
        x"6C41",
        x"206C",
        x"2000",
        x"6573",
        x"2074",
        x"7461",
        x"0020",
        x"7254",
        x"6361",
        x"6E69",
        x"2067",
        x"6964",
        x"6173",
        x"6C62",
        x"6465",
        x"000A",
        x"6920",
        x"736E",
        x"7274",
        x"6375",
        x"6974",
        x"6E6F",
        x"2073",
        x"6877",
        x"6C69",
        x"2065",
        x"6973",
        x"676E",
        x"656C",
        x"7320",
        x"6574",
        x"7070",
        x"6E69",
        x"0A67",
        x"5400",
        x"6172",
        x"6963",
        x"676E",
        x"6520",
        x"6576",
        x"7972",
        x"0020",
        x"7242",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"772F",
        x"7461",
        x"6863",
        x"6E20",
        x"746F",
        x"7320",
        x"7465",
        x"6120",
        x"2074",
        x"2000",
        x"6177",
        x"6374",
        x"6568",
        x"2F73",
        x"7262",
        x"6165",
        x"706B",
        x"696F",
        x"746E",
        x"2073",
        x"6D69",
        x"6C70",
        x"6D65",
        x"6E65",
        x"6574",
        x"0A64",
        x"4A00",
        x"6E75",
        x"3120",
        x"2037",
        x"3032",
        x"3032",
        x"2000",
        x"6E6F",
        x"0020",
        x"3731",
        x"323A",
        x"3A35",
        x"3935",
        x"0A00",
        x"6F43",
        x"706D",
        x"6C69",
        x"6465",
        x"6120",
        x"2074",
        x"3000",
        x"392E",
        x"3638",
        x"2000",
        x"6E49",
        x"432D",
        x"7269",
        x"7563",
        x"7469",
        x"4520",
        x"756D",
        x"616C",
        x"6F74",
        x"2072",
        x"6576",
        x"7372",
        x"6F69",
        x"206E",
        x"4900",
        x"4543",
        x"362D",
        x"4335",
        x"3230",
        x"2000",
        x"6572",
        x"6461",
        x"6E69",
        x"0067",
        x"7720",
        x"6972",
        x"6974",
        x"676E",
        x"2000",
        x"6968",
        x"2074",
        x"7461",
        x"0020",
        x"6420",
        x"6F72",
        x"7070",
        x"6465",
        x"000A",
        x"6520",
        x"6576",
        x"746E",
        x"3E00",
        x"003D",
        x"2020",
        x"2020",
        x"2020",
        x"2020",
        x"2020",
        x"203A",
        x"7400",
        x"6972",
        x"6767",
        x"7265",
        x"203A",
        x"4C49",
        x"454C",
        x"4147",
        x"004C",
        x"7274",
        x"6769",
        x"6567",
        x"3A72",
        x"0020",
        x"202C",
        x"2000",
        x"3E3C",
        x"0020",
        x"6E49",
        x"6F63",
        x"736E",
        x"7369",
        x"6574",
        x"746E",
        x"5220",
        x"3A64",
        x"0020",
        x"6452",
        x"203A",
        x"5700",
        x"3A72",
        x"0020",
        x"2020",
        x"5300",
        x"6E65",
        x"2064",
        x"6966",
        x"656C",
        x"6E20",
        x"776F",
        x"2E2E",
        x"0A2E",
        x"7500",
        x"6173",
        x"6567",
        x"0A3A",
        x"4900",
        x"6C6C",
        x"6765",
        x"6C61",
        x"6320",
        x"6D6F",
        x"616D",
        x"646E",
        x"203A",
        x"3E00",
        x"203E",
        x"9F00",
        x"3F82",
        x"A1BF",
        x"DF3F",
        x"3FC0",
        x"E0FF",
        x"E9F8",
        x"CBDA",
        x"ADBC",
        x"8F9E",
        x"6170",
        x"4352",
        x"2534",
        x"0716",
        x"B0A0",
        x"F0E0",
        x"9484",
        x"D4C4",
        x"3626",
        x"7666",
        x"1707",
        x"5747",
        x"9080",
        x"B0A0",
        x"D0C0",
        x"F0E0",
        x"1707",
        x"3727",
        x"5747",
        x"7767",
        x"D89C",
        x"9CF4",
        x"C488",
        x"4B88",
        x"283F",
        x"2433",
        x"021E",
        x"1C19",
        x"1293",
        x"1372",
        x"0028",
        x"0028",
        x"283F",
        x"2431",
        x"021E",
        x"1C19",
        x"0901",
        x"0967",
        x"000C",
        x"000C",
        x"283F",
        x"2431",
        x"0026",
        x"2320",
        x"0701",
        x"0867",
        x"000B",
        x"000B",
        x"507F",
        x"2862",
        x"021E",
        x"1C19",
        x"0901",
        x"0967",
        x"0008",
        x"0008",
        x"507F",
        x"2862",
        x"0026",
        x"2320",
        x"0701",
        x"0867",
        x"0006",
        x"0006",
        x"6C41",
        x"6177",
        x"7379",
        x"7E00",
        x"3054",
        x"6F20",
        x"2072",
        x"3154",
        x"5400",
        x"2030",
        x"6E78",
        x"726F",
        x"5420",
        x"0031",
        x"547E",
        x"2030",
        x"726F",
        x"7E20",
        x"3154",
        x"5400",
        x"2030",
        x"6F78",
        x"2072",
        x"3154",
        x"7E00",
        x"3054",
        x"7E00",
        x"3054",
        x"6120",
        x"646E",
        x"5420",
        x"0031",
        x"547E",
        x"2030",
        x"6E61",
        x"2064",
        x"547E",
        x"0031",
        x"654E",
        x"6576",
        x"0072",
        x"7254",
        x"6E61",
        x"6973",
        x"6E65",
        x"0074",
        x"7845",
        x"5720",
        x"7461",
        x"6863",
        x"4500",
        x"2078",
        x"7242",
        x"706B",
        x"0074",
        x"4F49",
        x"5720",
        x"2072",
        x"6157",
        x"6374",
        x"0068",
        x"4F49",
        x"5720",
        x"2072",
        x"7242",
        x"706B",
        x"0074",
        x"4F49",
        x"5220",
        x"2064",
        x"6157",
        x"6374",
        x"0068",
        x"4F49",
        x"5220",
        x"2064",
        x"7242",
        x"706B",
        x"0074",
        x"654D",
        x"206D",
        x"7257",
        x"5720",
        x"7461",
        x"6863",
        x"4D00",
        x"6D65",
        x"5720",
        x"2072",
        x"7242",
        x"706B",
        x"0074",
        x"654D",
        x"206D",
        x"6452",
        x"5720",
        x"7461",
        x"6863",
        x"4D00",
        x"6D65",
        x"5220",
        x"2064",
        x"7242",
        x"706B",
        x"0074",
        x"0712",
        x"0F11",
        x"0809",
        x"0118",
        x"0620",
        x"071B",
        x"0A0C",
        x"0710",
        x"0B0D",
        x"090B",
        x"0D0A",
        x"0D08",
        x"0116",
        x"021A",
        x"0329",
        x"000E",
        x"100F",
        x"0E17",
        x"0C21",
        x"0015",
        x"091D",
        x"071F",
        x"0E1E",
        x"071C",
        x"0622",
        x"0701",
        x"0406",
        x"0428",
        x"0404",
        x"0426",
        x"0405",
        x"0427",
        x"0007",
        x"0523",
        x"0000",
        x"07A5",
        x"0797",
        x"077D",
        x"0760",
        x"073D",
        x"0725",
        x"0712",
        x"0711",
        x"0705",
        x"06F7",
        x"06E1",
        x"06CC",
        x"06AF",
        x"069C",
        x"0690",
        x"0682",
        x"0668",
        x"6F3C",
        x"3170",
        x"203E",
        x"205B",
        x"6F3C",
        x"3270",
        x"203E",
        x"205B",
        x"6F3C",
        x"3370",
        x"203E",
        x"205D",
        x"005D",
        x"205B",
        x"633C",
        x"6D6F",
        x"616D",
        x"646E",
        x"203E",
        x"005D",
        x"205B",
        x"763C",
        x"6C61",
        x"6575",
        x"203E",
        x"005D",
        x"733C",
        x"6174",
        x"7472",
        x"203E",
        x"653C",
        x"646E",
        x"203E",
        x"743C",
        x"3E6F",
        x"3C00",
        x"7473",
        x"7261",
        x"3E74",
        x"3C20",
        x"6E65",
        x"3E64",
        x"5B20",
        x"3C20",
        x"6574",
        x"7473",
        x"6E20",
        x"6D75",
        x"203E",
        x"005D",
        x"733C",
        x"6174",
        x"7472",
        x"203E",
        x"653C",
        x"646E",
        x"203E",
        x"643C",
        x"7461",
        x"3E61",
        x"5B00",
        x"3C20",
        x"7473",
        x"7261",
        x"3E74",
        x"5B20",
        x"3C20",
        x"6E65",
        x"3E64",
        x"5D20",
        x"5D20",
        x"3C00",
        x"7473",
        x"7261",
        x"3E74",
        x"3C20",
        x"6E65",
        x"3E64",
        x"5B00",
        x"3C20",
        x"6572",
        x"6573",
        x"3E74",
        x"5D20",
        x"0000",
        x"205B",
        x"693C",
        x"736E",
        x"7274",
        x"6375",
        x"6974",
        x"6E6F",
        x"3E73",
        x"5D20",
        x"5B00",
        x"3C20",
        x"6461",
        x"7264",
        x"7365",
        x"3E73",
        x"3C20",
        x"7274",
        x"6769",
        x"6567",
        x"3E72",
        x"5D20",
        x"3C00",
        x"6461",
        x"7264",
        x"7365",
        x"3E73",
        x"5B20",
        x"3C20",
        x"616D",
        x"6B73",
        x"203E",
        x"205B",
        x"743C",
        x"6972",
        x"6767",
        x"7265",
        x"203E",
        x"205D",
        x"005D",
        x"613C",
        x"6464",
        x"6572",
        x"7373",
        x"203E",
        x"643C",
        x"7461",
        x"3E61",
        x"5B20",
        x"3C20",
        x"6F63",
        x"6E75",
        x"3E74",
        x"5D20",
        x"5B00",
        x"3C20",
        x"6461",
        x"7264",
        x"7365",
        x"3E73",
        x"5B20",
        x"3C20",
        x"6F63",
        x"6E75",
        x"3E74",
        x"5D20",
        x"5D20",
        x"5B00",
        x"3C20",
        x"6461",
        x"7264",
        x"7365",
        x"3E73",
        x"5D20",
        x"3C00",
        x"6461",
        x"7264",
        x"7365",
        x"3E73",
        x"0000",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"010E",
        x"0C00",
        x"0D0D",
        x"0C00",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0606",
        x"0000",
        x"010E",
        x"0D00",
        x"0D0D",
        x"0000",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0000",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0104",
        x"0F00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0606",
        x"0000",
        x"000E",
        x"1000",
        x"0D0D",
        x"0300",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0706",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0400",
        x"0408",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0600",
        x"0706",
        x"0000",
        x"000E",
        x"0D00",
        x"0E0D",
        x"0400",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0400",
        x"0008",
        x"0500",
        x"0505",
        x"0000",
        x"0004",
        x"0C00",
        x"0C0C",
        x"0300",
        x"0A09",
        x"0500",
        x"0606",
        x"0000",
        x"000E",
        x"0C00",
        x"0D0D",
        x"0B00",
        x"4223",
        x"3C42",
        x"0223",
        x"2542",
        x"0223",
        x"3C42",
        x"0223",
        x"0942",
        x"2323",
        x"3B42",
        x"0223",
        x"0E42",
        x"1923",
        x"3B42",
        x"0223",
        x"1D42",
        x"4201",
        x"0642",
        x"2C01",
        x"2942",
        x"2C01",
        x"0642",
        x"2C01",
        x"0742",
        x"0101",
        x"0642",
        x"2C01",
        x"3142",
        x"1501",
        x"0642",
        x"2C01",
        x"2E42",
        x"4218",
        x"4242",
        x"2118",
        x"2442",
        x"2118",
        x"1C42",
        x"2118",
        x"0C42",
        x"1818",
        x"4242",
        x"2118",
        x"1042",
        x"2718",
        x"4242",
        x"2118",
        x"2F42",
        x"4200",
        x"3842",
        x"2D00",
        x"2842",
        x"2D00",
        x"1C42",
        x"2D00",
        x"0D42",
        x"0000",
        x"3842",
        x"2D00",
        x"3342",
        x"2B00",
        x"1C42",
        x"2D00",
        x"0A42",
        x"4234",
        x"3742",
        x"3634",
        x"1742",
        x"3E06",
        x"3742",
        x"3634",
        x"0342",
        x"3434",
        x"3742",
        x"3634",
        x"4042",
        x"3F34",
        x"3842",
        x"3834",
        x"2042",
        x"1F1E",
        x"2042",
        x"1F1E",
        x"3A42",
        x"391E",
        x"2042",
        x"1F1E",
        x"0442",
        x"1E1E",
        x"2042",
        x"1F1E",
        x"1142",
        x"3D1E",
        x"2042",
        x"1F1E",
        x"1442",
        x"4212",
        x"1442",
        x"1512",
        x"1B42",
        x"1612",
        x"1441",
        x"1512",
        x"0842",
        x"1212",
        x"4242",
        x"1512",
        x"0F42",
        x"2612",
        x"4235",
        x"1512",
        x"1342",
        x"4230",
        x"1342",
        x"1930",
        x"1A42",
        x"2230",
        x"1342",
        x"1930",
        x"0542",
        x"3030",
        x"4242",
        x"1930",
        x"3242",
        x"2A30",
        x"4242",
        x"1930",
        x"4142",
        x"4344",
        x"4E41",
        x"4144",
        x"4C53",
        x"4342",
        x"4243",
        x"5343",
        x"4542",
        x"4251",
        x"5449",
        x"4D42",
        x"4249",
        x"454E",
        x"5042",
        x"424C",
        x"4152",
        x"5242",
        x"424B",
        x"4356",
        x"5642",
        x"4353",
        x"434C",
        x"4C43",
        x"4344",
        x"494C",
        x"4C43",
        x"4356",
        x"504D",
        x"5043",
        x"4358",
        x"5950",
        x"4544",
        x"4443",
        x"5845",
        x"4544",
        x"4559",
        x"524F",
        x"4E49",
        x"4943",
        x"584E",
        x"4E49",
        x"4A59",
        x"504D",
        x"534A",
        x"4C52",
        x"4144",
        x"444C",
        x"4C58",
        x"5944",
        x"534C",
        x"4E52",
        x"504F",
        x"524F",
        x"5041",
        x"4148",
        x"4850",
        x"5050",
        x"5848",
        x"4850",
        x"5059",
        x"414C",
        x"4C50",
        x"5050",
        x"584C",
        x"4C50",
        x"5259",
        x"4C4F",
        x"4F52",
        x"5252",
        x"4954",
        x"5452",
        x"5353",
        x"4342",
        x"4553",
        x"5343",
        x"4445",
        x"4553",
        x"5349",
        x"4154",
        x"5453",
        x"5350",
        x"5854",
        x"5453",
        x"5359",
        x"5A54",
        x"4154",
        x"5458",
        x"5941",
        x"5254",
        x"5442",
        x"4253",
        x"5354",
        x"5458",
        x"4158",
        x"5854",
        x"5453",
        x"4159",
        x"4157",
        x"2D49",
        x"2D2D",
        x"2000",
        x"5320",
        x"6174",
        x"7574",
        x"3A73",
        x"0020",
        x"5020",
        x"3D43",
        x"2000",
        x"5053",
        x"303D",
        x"0031",
        x"5920",
        x"003D",
        x"5820",
        x"003D",
        x"3536",
        x"3230",
        x"5220",
        x"6765",
        x"7369",
        x"6574",
        x"7372",
        x"0A3A",
        x"2020",
        x"3D41",
        x"0000",
        x"2411",
        x"BE1F",
        x"EFCF",
        x"E0DF",
        x"BFDE",
        x"BFCD",
        x"E012",
        x"E6A0",
        x"E0B0",
        x"E2E2",
        x"E3F8",
        x"EF0F",
        x"9503",
        x"BF0B",
        x"C004",
        x"95D8",
        x"920D",
        x"9631",
        x"F3C8",
        x"39A4",
        x"07B1",
        x"F7C9",
        x"E024",
        x"E9A4",
        x"E0B2",
        x"C001",
        x"921D",
        x"3FA8",
        x"07B2",
        x"F7E1",
        x"940E",
        x"19E5",
        x"940C",
        x"1C0F",
        x"940C",
        x"0000",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"E001",
        x"E010",
        x"24FF",
        x"94F3",
        x"9180",
        x"0060",
        x"2FC0",
        x"2FD1",
        x"0FC8",
        x"1DD1",
        x"FD87",
        x"95DA",
        x"70CF",
        x"27DD",
        x"E085",
        x"0FCC",
        x"1FDD",
        x"958A",
        x"F7E1",
        x"54C5",
        x"4FDD",
        x"8188",
        x"2388",
        x"F0B1",
        x"E58B",
        x"940E",
        x"162A",
        x"24EE",
        x"94E3",
        x"0CEF",
        x"2D8F",
        x"E090",
        x"940E",
        x"16C0",
        x"E880",
        x"E090",
        x"940E",
        x"1652",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"162D",
        x"E08A",
        x"940E",
        x"162A",
        x"2CFE",
        x"5F0F",
        x"4F1F",
        x"3101",
        x"0511",
        x"F689",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"1AE9",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2EE8",
        x"2EF9",
        x"2FC6",
        x"E08D",
        x"940E",
        x"160F",
        x"E18B",
        x"940E",
        x"160F",
        x"E58B",
        x"940E",
        x"160F",
        x"E48B",
        x"940E",
        x"160F",
        x"E987",
        x"E094",
        x"940E",
        x"1652",
        x"23CC",
        x"F081",
        x"2D0E",
        x"2D1F",
        x"2FC0",
        x"2FD1",
        x"19CE",
        x"09DF",
        x"2FE0",
        x"2FF1",
        x"9181",
        x"2F0E",
        x"2F1F",
        x"2388",
        x"F029",
        x"940E",
        x"160F",
        x"CFF2",
        x"E0C0",
        x"E0D0",
        x"E000",
        x"940E",
        x"1623",
        x"2F18",
        x"3002",
        x"F439",
        x"3481",
        x"F409",
        x"C03F",
        x"3482",
        x"F7A9",
        x"E081",
        x"C03C",
        x"3001",
        x"F421",
        x"358B",
        x"F779",
        x"E002",
        x"CFEE",
        x"318B",
        x"F411",
        x"5F0F",
        x"CFEA",
        x"3088",
        x"F469",
        x"9720",
        x"F331",
        x"9721",
        x"E088",
        x"940E",
        x"160F",
        x"E280",
        x"940E",
        x"160F",
        x"E088",
        x"940E",
        x"160F",
        x"CFDB",
        x"308D",
        x"F4A9",
        x"9720",
        x"F441",
        x"2DCE",
        x"2DDF",
        x"9189",
        x"2388",
        x"F031",
        x"940E",
        x"160F",
        x"CFFA",
        x"0DCE",
        x"1DDF",
        x"8218",
        x"E08A",
        x"940E",
        x"160F",
        x"E08D",
        x"940E",
        x"160F",
        x"E080",
        x"C00C",
        x"3280",
        x"F214",
        x"940E",
        x"160F",
        x"2DEE",
        x"2DFF",
        x"0FEC",
        x"1FFD",
        x"8310",
        x"9621",
        x"CFB9",
        x"EF8F",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"1AE9",
        x"E0A0",
        x"E0B0",
        x"E3EA",
        x"E0F6",
        x"940C",
        x"1AC9",
        x"2EC8",
        x"2ED9",
        x"2FA8",
        x"2FB9",
        x"910D",
        x"911C",
        x"2CA1",
        x"2FC0",
        x"2FD1",
        x"0DCA",
        x"1DD1",
        x"8188",
        x"5681",
        x"318A",
        x"F410",
        x"94A3",
        x"CFF6",
        x"EB82",
        x"2EE8",
        x"E080",
        x"2EF8",
        x"2CB1",
        x"2DEE",
        x"2DFF",
        x"9181",
        x"9191",
        x"2EEE",
        x"2EFF",
        x"2FE8",
        x"2FF9",
        x"9001",
        x"2000",
        x"F7E9",
        x"9731",
        x"1BE8",
        x"16AE",
        x"F408",
        x"2DEA",
        x"2F4E",
        x"E050",
        x"2F60",
        x"2F71",
        x"940E",
        x"1B74",
        x"2B89",
        x"F461",
        x"2FEC",
        x"2FFD",
        x"9621",
        x"8180",
        x"3280",
        x"F3D1",
        x"2DAC",
        x"2DBD",
        x"93ED",
        x"93FC",
        x"2D8B",
        x"C005",
        x"94B3",
        x"E2B2",
        x"16BB",
        x"F6C1",
        x"EF8F",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"1AE5",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"E885",
        x"E094",
        x"940E",
        x"1652",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"162D",
        x"E08A",
        x"940E",
        x"162A",
        x"91DF",
        x"91CF",
        x"9508",
        x"B330",
        x"2B86",
        x"2B97",
        x"B328",
        x"7E20",
        x"BB28",
        x"B328",
        x"2F48",
        x"6240",
        x"2724",
        x"BB28",
        x"E140",
        x"E257",
        x"5041",
        x"0951",
        x"F029",
        x"B320",
        x"2723",
        x"FF26",
        x"CFF9",
        x"9508",
        x"9190",
        x"0294",
        x"FF84",
        x"C002",
        x"6092",
        x"C001",
        x"6091",
        x"9390",
        x"0294",
        x"9508",
        x"E060",
        x"E070",
        x"E182",
        x"E090",
        x"940E",
        x"0690",
        x"9508",
        x"EF80",
        x"E091",
        x"940E",
        x"1652",
        x"E060",
        x"E070",
        x"E08A",
        x"E090",
        x"940E",
        x"0690",
        x"9508",
        x"B392",
        x"7C90",
        x"BB92",
        x"B392",
        x"2B89",
        x"BB82",
        x"E088",
        x"958A",
        x"F7F1",
        x"B181",
        x"9508",
        x"E060",
        x"E070",
        x"E180",
        x"E090",
        x"940E",
        x"0690",
        x"E082",
        x"940E",
        x"06C1",
        x"9508",
        x"E060",
        x"E070",
        x"E181",
        x"E090",
        x"940E",
        x"0690",
        x"E082",
        x"940E",
        x"06C1",
        x"9508",
        x"B392",
        x"7C90",
        x"BB92",
        x"B392",
        x"2B89",
        x"BB82",
        x"E088",
        x"958A",
        x"F7F1",
        x"B181",
        x"9A90",
        x"E098",
        x"959A",
        x"F7F1",
        x"B121",
        x"E090",
        x"2B92",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"2F08",
        x"2F19",
        x"2FC6",
        x"23CC",
        x"F061",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E084",
        x"E090",
        x"940E",
        x"0690",
        x"9516",
        x"9507",
        x"50C1",
        x"CFF2",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"2EE6",
        x"2EF7",
        x"2F04",
        x"2F15",
        x"2FC2",
        x"E160",
        x"940E",
        x"06F2",
        x"E160",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"06F2",
        x"E06A",
        x"2F80",
        x"2F91",
        x"940E",
        x"06F2",
        x"E064",
        x"2F8C",
        x"E090",
        x"940E",
        x"06F2",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"9508",
        x"E68B",
        x"E094",
        x"940E",
        x"1652",
        x"9508",
        x"EE90",
        x"0F98",
        x"359F",
        x"F008",
        x"E28E",
        x"940E",
        x"162A",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"2F08",
        x"2F19",
        x"2FC6",
        x"E280",
        x"940E",
        x"162A",
        x"2F80",
        x"2F91",
        x"940E",
        x"167A",
        x"E38A",
        x"940E",
        x"162A",
        x"2F8C",
        x"940E",
        x"166F",
        x"E688",
        x"E094",
        x"940E",
        x"1652",
        x"2F8C",
        x"940E",
        x"0731",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FD8",
        x"E0C8",
        x"2F6D",
        x"7061",
        x"E070",
        x"E08C",
        x"E090",
        x"940E",
        x"0690",
        x"95D6",
        x"50C1",
        x"F7B1",
        x"91DF",
        x"91CF",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"2F08",
        x"2F19",
        x"E1C0",
        x"2F60",
        x"2F71",
        x"7061",
        x"2777",
        x"E08C",
        x"E090",
        x"940E",
        x"0690",
        x"9516",
        x"9507",
        x"50C1",
        x"F7A1",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"E8E4",
        x"E0F7",
        x"940C",
        x"1AD0",
        x"9120",
        x"0297",
        x"9130",
        x"0298",
        x"833C",
        x"832B",
        x"821A",
        x"8219",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"17D9",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17D9",
        x"818B",
        x"819C",
        x"9390",
        x"0298",
        x"9380",
        x"0297",
        x"940E",
        x"0768",
        x"E010",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"1821",
        x"9390",
        x"0298",
        x"9380",
        x"0297",
        x"5F1F",
        x"8129",
        x"813A",
        x"1521",
        x"0531",
        x"F419",
        x"301A",
        x"F370",
        x"C008",
        x"814B",
        x"815C",
        x"1748",
        x"0759",
        x"F418",
        x"1728",
        x"0739",
        x"F728",
        x"9624",
        x"E0E3",
        x"940C",
        x"1AEC",
        x"E060",
        x"E070",
        x"E183",
        x"E090",
        x"940E",
        x"0690",
        x"9508",
        x"E060",
        x"E070",
        x"E184",
        x"E090",
        x"940E",
        x"0690",
        x"E082",
        x"940E",
        x"06C1",
        x"9508",
        x"E060",
        x"E070",
        x"E185",
        x"E090",
        x"940E",
        x"0690",
        x"E082",
        x"940E",
        x"06C1",
        x"9508",
        x"E060",
        x"E070",
        x"E186",
        x"E090",
        x"940E",
        x"0690",
        x"9508",
        x"E060",
        x"E070",
        x"E187",
        x"E090",
        x"940E",
        x"0690",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"940E",
        x"0768",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1821",
        x"91DF",
        x"91CF",
        x"9508",
        x"E1A0",
        x"E0B0",
        x"EFEC",
        x"E0F7",
        x"940C",
        x"1AC7",
        x"2E86",
        x"2E97",
        x"E967",
        x"E072",
        x"940E",
        x"17D9",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"0768",
        x"2CE1",
        x"2CF1",
        x"2EAC",
        x"2EBD",
        x"E181",
        x"0EA8",
        x"1CB1",
        x"2F0C",
        x"2F1D",
        x"5F0F",
        x"4F1F",
        x"2EC0",
        x"2ED1",
        x"2DE8",
        x"2DF9",
        x"9509",
        x"2DEC",
        x"2DFD",
        x"9381",
        x"2ECE",
        x"2EDF",
        x"15EA",
        x"05FB",
        x"F7A9",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"0D8E",
        x"1D9F",
        x"940E",
        x"167A",
        x"E280",
        x"940E",
        x"162A",
        x"2EC0",
        x"2ED1",
        x"2DEC",
        x"2DFD",
        x"9181",
        x"2ECE",
        x"2EDF",
        x"940E",
        x"166F",
        x"E280",
        x"940E",
        x"162A",
        x"14CA",
        x"04DB",
        x"F799",
        x"E280",
        x"940E",
        x"162A",
        x"2FE0",
        x"2FF1",
        x"9181",
        x"2F0E",
        x"2F1F",
        x"940E",
        x"0731",
        x"150A",
        x"051B",
        x"F7B1",
        x"E08A",
        x"940E",
        x"162A",
        x"E1F0",
        x"0EEF",
        x"1CF1",
        x"14E1",
        x"E081",
        x"06F8",
        x"F009",
        x"CFBD",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"9593",
        x"9390",
        x"0298",
        x"9380",
        x"0297",
        x"9660",
        x"E0EC",
        x"940C",
        x"1AE3",
        x"ED66",
        x"E076",
        x"940E",
        x"07F6",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"E6EA",
        x"E0F8",
        x"940C",
        x"1ACA",
        x"2EE6",
        x"2EF7",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"E967",
        x"E072",
        x"940E",
        x"17D9",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"1768",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"0768",
        x"2DEE",
        x"2DFF",
        x"9509",
        x"2ED8",
        x"2F08",
        x"E010",
        x"E58E",
        x"E094",
        x"940E",
        x"1652",
        x"2D6D",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"0739",
        x"E08A",
        x"940E",
        x"162A",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"5041",
        x"0951",
        x"0961",
        x"0971",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"9702",
        x"05A1",
        x"05B1",
        x"F0EC",
        x"2DEE",
        x"2DFF",
        x"9509",
        x"2EB8",
        x"2EC8",
        x"2CD1",
        x"150C",
        x"051D",
        x"F089",
        x"E48C",
        x"E094",
        x"940E",
        x"1652",
        x"2D8B",
        x"940E",
        x"166F",
        x"E487",
        x"E094",
        x"940E",
        x"1652",
        x"2F80",
        x"940E",
        x"166F",
        x"E08A",
        x"940E",
        x"162A",
        x"2D0C",
        x"2D1D",
        x"CFCF",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"9601",
        x"9390",
        x"0298",
        x"9380",
        x"0297",
        x"9624",
        x"E0E9",
        x"940C",
        x"1AE6",
        x"EC6C",
        x"E076",
        x"940E",
        x"0864",
        x"9508",
        x"E1A0",
        x"E0B0",
        x"EEE1",
        x"E0F8",
        x"940C",
        x"1ACB",
        x"2F08",
        x"2F86",
        x"940E",
        x"06C1",
        x"2F18",
        x"2F80",
        x"940E",
        x"06E0",
        x"2F48",
        x"2F59",
        x"E060",
        x"E070",
        x"2B61",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"2EE8",
        x"2EF9",
        x"940E",
        x"16D6",
        x"2DEE",
        x"2DFF",
        x"9001",
        x"2000",
        x"F7E9",
        x"9731",
        x"19EE",
        x"09FF",
        x"E000",
        x"E010",
        x"E088",
        x"E090",
        x"2EC8",
        x"2ED9",
        x"1ACE",
        x"08D1",
        x"150C",
        x"051D",
        x"F414",
        x"E380",
        x"C007",
        x"2FE0",
        x"2FF1",
        x"19EC",
        x"09FD",
        x"0DEE",
        x"1DFF",
        x"8180",
        x"940E",
        x"162A",
        x"3007",
        x"0511",
        x"F041",
        x"3001",
        x"F419",
        x"E28E",
        x"940E",
        x"162A",
        x"5F0F",
        x"4F1F",
        x"CFE7",
        x"E682",
        x"E091",
        x"940E",
        x"162D",
        x"9660",
        x"E0E8",
        x"940C",
        x"1AE7",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2F08",
        x"2F19",
        x"E4CC",
        x"E0D1",
        x"E622",
        x"2EE2",
        x"E021",
        x"2EF2",
        x"E081",
        x"FF00",
        x"C00B",
        x"2388",
        x"F421",
        x"E484",
        x"E094",
        x"940E",
        x"1652",
        x"8188",
        x"8199",
        x"940E",
        x"1652",
        x"E080",
        x"9516",
        x"9507",
        x"9622",
        x"16EC",
        x"06FD",
        x"F769",
        x"B7CD",
        x"B7DE",
        x"E0E6",
        x"940C",
        x"1AE9",
        x"93CF",
        x"2FC8",
        x"3180",
        x"F468",
        x"E38A",
        x"E094",
        x"940E",
        x"1652",
        x"2FEC",
        x"E0F0",
        x"0FEE",
        x"1FFF",
        x"5DE4",
        x"4FFE",
        x"8180",
        x"8191",
        x"C002",
        x"E289",
        x"E094",
        x"940E",
        x"1652",
        x"91CF",
        x"9508",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"9180",
        x"0299",
        x"9190",
        x"029A",
        x"2B89",
        x"F409",
        x"C046",
        x"2CF1",
        x"2DCF",
        x"E0D0",
        x"9180",
        x"0299",
        x"9190",
        x"029A",
        x"17C8",
        x"07D9",
        x"F00C",
        x"C03F",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"16C0",
        x"E186",
        x"E091",
        x"940E",
        x"1652",
        x"2F0C",
        x"2F1D",
        x"0F00",
        x"1F11",
        x"2FE0",
        x"2FF1",
        x"52E8",
        x"4FFB",
        x"8180",
        x"8191",
        x"940E",
        x"167A",
        x"E08F",
        x"E091",
        x"940E",
        x"1652",
        x"2FE0",
        x"2FF1",
        x"53E9",
        x"4FFB",
        x"8180",
        x"8191",
        x"940E",
        x"167A",
        x"E08C",
        x"E091",
        x"940E",
        x"1652",
        x"2FE0",
        x"2FF1",
        x"51E8",
        x"4FFB",
        x"8180",
        x"8191",
        x"940E",
        x"0926",
        x"E686",
        x"E091",
        x"940E",
        x"162D",
        x"54C5",
        x"4FDB",
        x"8188",
        x"940E",
        x"094D",
        x"E089",
        x"E091",
        x"940E",
        x"1652",
        x"94F3",
        x"CFBB",
        x"EF85",
        x"E090",
        x"940E",
        x"1652",
        x"B7CD",
        x"B7DE",
        x"E0E5",
        x"940C",
        x"1AEA",
        x"E0A0",
        x"E0B0",
        x"ECE5",
        x"E0F9",
        x"940C",
        x"1AC9",
        x"E086",
        x"940E",
        x"06E0",
        x"2EE8",
        x"2EF9",
        x"E088",
        x"940E",
        x"06E0",
        x"2EC8",
        x"2ED9",
        x"E08A",
        x"940E",
        x"06C1",
        x"2EA8",
        x"E08B",
        x"940E",
        x"06C1",
        x"2FC8",
        x"7081",
        x"2EB8",
        x"2F0C",
        x"E010",
        x"E084",
        x"9516",
        x"9507",
        x"958A",
        x"F7E1",
        x"2FD0",
        x"2300",
        x"F0D9",
        x"E18C",
        x"E094",
        x"940E",
        x"1652",
        x"300F",
        x"F421",
        x"E189",
        x"E094",
        x"940E",
        x"1652",
        x"2F80",
        x"2F91",
        x"940E",
        x"16C0",
        x"E182",
        x"E094",
        x"940E",
        x"1652",
        x"30D1",
        x"F019",
        x"E783",
        x"940E",
        x"162A",
        x"E088",
        x"E094",
        x"940E",
        x"1652",
        x"2F8C",
        x"708F",
        x"E0C1",
        x"E0D0",
        x"C002",
        x"0FCC",
        x"1FDD",
        x"958A",
        x"F7E2",
        x"2F8C",
        x"2F9D",
        x"7A8A",
        x"7092",
        x"2B89",
        x"F031",
        x"E06E",
        x"E070",
        x"E08C",
        x"E090",
        x"940E",
        x"08DB",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"0926",
        x"EF8F",
        x"E093",
        x"940E",
        x"1652",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"167A",
        x"23CC",
        x"F091",
        x"2F8C",
        x"2F9D",
        x"7C8C",
        x"2799",
        x"2B89",
        x"F019",
        x"EF86",
        x"E093",
        x"C002",
        x"EE8D",
        x"E093",
        x"940E",
        x"1652",
        x"2D6A",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"0739",
        x"E08A",
        x"940E",
        x"162A",
        x"75C5",
        x"27DD",
        x"2BCD",
        x"F051",
        x"E06E",
        x"E070",
        x"E08C",
        x"E090",
        x"940E",
        x"08DB",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"07E9",
        x"2D8B",
        x"B7CD",
        x"B7DE",
        x"E0EA",
        x"940C",
        x"1AE5",
        x"E587",
        x"E092",
        x"9701",
        x"F7F1",
        x"C000",
        x"0000",
        x"E080",
        x"940E",
        x"06E0",
        x"9390",
        x"0298",
        x"9380",
        x"0297",
        x"E063",
        x"E070",
        x"E084",
        x"E090",
        x"940E",
        x"08DB",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"07E9",
        x"9390",
        x"0296",
        x"9380",
        x"0295",
        x"9508",
        x"EE83",
        x"E093",
        x"940E",
        x"1652",
        x"EC85",
        x"E093",
        x"940E",
        x"1652",
        x"EB8F",
        x"E093",
        x"940E",
        x"1652",
        x"EB81",
        x"E093",
        x"940E",
        x"1652",
        x"EA88",
        x"E093",
        x"940E",
        x"1652",
        x"EA83",
        x"E093",
        x"940E",
        x"1652",
        x"E987",
        x"E093",
        x"940E",
        x"1652",
        x"E08A",
        x"940E",
        x"162A",
        x"E088",
        x"E090",
        x"940E",
        x"16C0",
        x"E785",
        x"E093",
        x"940E",
        x"1652",
        x"9508",
        x"9140",
        x"0299",
        x"9150",
        x"029A",
        x"EDE8",
        x"E0F4",
        x"E020",
        x"E030",
        x"1724",
        x"0735",
        x"F45C",
        x"9161",
        x"9171",
        x"1786",
        x"0797",
        x"F419",
        x"2F82",
        x"2F93",
        x"C003",
        x"5F2F",
        x"4F3F",
        x"CFF2",
        x"1784",
        x"0795",
        x"F010",
        x"EF8F",
        x"EF9F",
        x"9508",
        x"E061",
        x"E070",
        x"2388",
        x"F411",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"0690",
        x"9508",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"1616",
        x"0617",
        x"0618",
        x"0619",
        x"F47C",
        x"E489",
        x"E093",
        x"940E",
        x"1652",
        x"2D9F",
        x"2D8E",
        x"2D7D",
        x"2D6C",
        x"940E",
        x"16E2",
        x"E284",
        x"E093",
        x"940E",
        x"1652",
        x"C008",
        x"E182",
        x"E093",
        x"940E",
        x"1652",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"92C0",
        x"04C3",
        x"92D0",
        x"04C4",
        x"92E0",
        x"04C5",
        x"92F0",
        x"04C6",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"9508",
        x"E0A4",
        x"E0B0",
        x"EEEE",
        x"E0FA",
        x"940C",
        x"1AD1",
        x"9140",
        x"04C3",
        x"9150",
        x"04C4",
        x"9160",
        x"04C5",
        x"9170",
        x"04C6",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"1768",
        x"8169",
        x"817A",
        x"818B",
        x"819C",
        x"940E",
        x"0AB7",
        x"9624",
        x"E0E2",
        x"940C",
        x"1AED",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F86",
        x"2F97",
        x"940E",
        x"0926",
        x"E089",
        x"E093",
        x"940E",
        x"1652",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"91DF",
        x"91CF",
        x"9508",
        x"E084",
        x"E093",
        x"940E",
        x"1652",
        x"9180",
        x"0299",
        x"9190",
        x"029A",
        x"940E",
        x"16C0",
        x"EE86",
        x"E092",
        x"940E",
        x"1652",
        x"9508",
        x"93CF",
        x"E060",
        x"E070",
        x"E082",
        x"E090",
        x"940E",
        x"0690",
        x"E0C0",
        x"2F8C",
        x"E090",
        x"9120",
        x"0299",
        x"9130",
        x"029A",
        x"1782",
        x"0793",
        x"F4EC",
        x"2FE8",
        x"2FF9",
        x"54E5",
        x"4FFB",
        x"0F88",
        x"1F99",
        x"2FA8",
        x"2FB9",
        x"51A8",
        x"4FBB",
        x"914D",
        x"915C",
        x"2FA8",
        x"2FB9",
        x"53A9",
        x"4FBB",
        x"916D",
        x"917C",
        x"2FA8",
        x"2FB9",
        x"52A8",
        x"4FBB",
        x"8120",
        x"918D",
        x"919C",
        x"940E",
        x"070A",
        x"5FCF",
        x"CFDA",
        x"2FC2",
        x"30C8",
        x"F458",
        x"E020",
        x"E040",
        x"E050",
        x"E060",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"070A",
        x"5FCF",
        x"CFF3",
        x"E061",
        x"E070",
        x"E082",
        x"E090",
        x"940E",
        x"0690",
        x"91CF",
        x"9508",
        x"930F",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"2FAE",
        x"2FBF",
        x"52A8",
        x"4FBB",
        x"2364",
        x"2375",
        x"936D",
        x"937C",
        x"2FAE",
        x"2FBF",
        x"53A9",
        x"4FBB",
        x"934D",
        x"935C",
        x"51E8",
        x"4FFB",
        x"8331",
        x"8320",
        x"2FE8",
        x"2FF9",
        x"54E5",
        x"4FFB",
        x"8300",
        x"940E",
        x"0B2F",
        x"910F",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"9120",
        x"0299",
        x"9130",
        x"029A",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"2FAE",
        x"2FBF",
        x"52A8",
        x"4FBB",
        x"2FCE",
        x"2FDF",
        x"53C9",
        x"4FDB",
        x"2F0E",
        x"2F1F",
        x"5108",
        x"4F1B",
        x"2F48",
        x"2F59",
        x"5445",
        x"4F5B",
        x"1782",
        x"0793",
        x"F4D4",
        x"9601",
        x"9612",
        x"916D",
        x"917C",
        x"9713",
        x"936D",
        x"937D",
        x"816A",
        x"817B",
        x"9369",
        x"9379",
        x"2FE0",
        x"2FF1",
        x"8162",
        x"8173",
        x"9361",
        x"9371",
        x"2F0E",
        x"2F1F",
        x"2FE4",
        x"2FF5",
        x"8161",
        x"9361",
        x"2F4E",
        x"2F5F",
        x"CFE3",
        x"5021",
        x"0931",
        x"9330",
        x"029A",
        x"9320",
        x"0299",
        x"940E",
        x"0B2F",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"3F6F",
        x"EF2F",
        x"0772",
        x"F419",
        x"FF80",
        x"C01D",
        x"C01E",
        x"3F6E",
        x"EF2F",
        x"0772",
        x"F419",
        x"FF80",
        x"C018",
        x"C015",
        x"3F6D",
        x"EF2F",
        x"0772",
        x"F411",
        x"EC63",
        x"C005",
        x"3F6C",
        x"EF2F",
        x"0772",
        x"F421",
        x"E36C",
        x"2786",
        x"2789",
        x"9508",
        x"FF77",
        x"C003",
        x"940E",
        x"1B50",
        x"9508",
        x"2F86",
        x"9508",
        x"EA8A",
        x"9508",
        x"E585",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E0E6",
        x"E0FC",
        x"940C",
        x"1AC1",
        x"2E28",
        x"2E39",
        x"2F06",
        x"2F17",
        x"2FC4",
        x"2FD5",
        x"2F84",
        x"2F95",
        x"940E",
        x"1B55",
        x"2CC2",
        x"2CD3",
        x"2CE1",
        x"2CF1",
        x"2C8C",
        x"2C9D",
        x"2CAE",
        x"2CBF",
        x"2E40",
        x"2E51",
        x"2C61",
        x"2C71",
        x"1448",
        x"0459",
        x"046A",
        x"047B",
        x"F0A4",
        x"2F6C",
        x"2F7D",
        x"2D88",
        x"2D99",
        x"940E",
        x"0BD9",
        x"940E",
        x"0757",
        x"2D88",
        x"2D99",
        x"940E",
        x"0768",
        x"940E",
        x"07C0",
        x"EF8F",
        x"1A88",
        x"0A98",
        x"0AA8",
        x"0AB8",
        x"CFE7",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"1B55",
        x"2D82",
        x"2D93",
        x"940E",
        x"0768",
        x"E000",
        x"E010",
        x"144C",
        x"045D",
        x"046E",
        x"047F",
        x"F174",
        x"940E",
        x"06D6",
        x"2EB8",
        x"2F6C",
        x"2F7D",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"0BD9",
        x"2EA8",
        x"16B8",
        x"F0E1",
        x"EC8C",
        x"E092",
        x"940E",
        x"1652",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"167A",
        x"EC82",
        x"E092",
        x"940E",
        x"1652",
        x"2D8A",
        x"940E",
        x"166F",
        x"EB85",
        x"E092",
        x"940E",
        x"1652",
        x"2D8B",
        x"940E",
        x"166F",
        x"EB82",
        x"E092",
        x"940E",
        x"1652",
        x"5F0F",
        x"4F1F",
        x"EF8F",
        x"1AC8",
        x"0AD8",
        x"0AE8",
        x"0AF8",
        x"CFCD",
        x"24EE",
        x"24FF",
        x"1AEC",
        x"0AFD",
        x"FCF7",
        x"C008",
        x"E086",
        x"16E8",
        x"04F1",
        x"F034",
        x"E095",
        x"2EE9",
        x"2CF1",
        x"C002",
        x"2CE1",
        x"2CF1",
        x"EA84",
        x"E092",
        x"940E",
        x"1652",
        x"2DEE",
        x"2DFF",
        x"0FEE",
        x"1FFF",
        x"59EF",
        x"4FFF",
        x"8180",
        x"8191",
        x"940E",
        x"162D",
        x"FDD7",
        x"C006",
        x"E280",
        x"940E",
        x"162A",
        x"2F8C",
        x"940E",
        x"166F",
        x"1501",
        x"0511",
        x"F059",
        x"E989",
        x"E092",
        x"940E",
        x"1652",
        x"2F80",
        x"2F91",
        x"940E",
        x"16C0",
        x"E980",
        x"E092",
        x"C002",
        x"E886",
        x"E092",
        x"940E",
        x"1652",
        x"B7CD",
        x"B7DE",
        x"E1E2",
        x"940C",
        x"1ADD",
        x"93CF",
        x"9B87",
        x"C00A",
        x"940E",
        x"09BF",
        x"2FC8",
        x"E060",
        x"E070",
        x"E089",
        x"E090",
        x"940E",
        x"0690",
        x"C001",
        x"E0C1",
        x"940E",
        x"1627",
        x"2388",
        x"F029",
        x"940E",
        x"1623",
        x"308D",
        x"F409",
        x"E0C0",
        x"2F8C",
        x"91CF",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"1768",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"1618",
        x"0619",
        x"061A",
        x"061B",
        x"F02C",
        x"E480",
        x"E092",
        x"940E",
        x"1652",
        x"C06C",
        x"E386",
        x"E092",
        x"940E",
        x"1652",
        x"8169",
        x"817A",
        x"818B",
        x"819C",
        x"940E",
        x"16E2",
        x"E287",
        x"E092",
        x"940E",
        x"1652",
        x"9080",
        x"04C3",
        x"9090",
        x"04C4",
        x"90A0",
        x"04C5",
        x"90B0",
        x"04C6",
        x"24CC",
        x"94C3",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F40C",
        x"C047",
        x"E060",
        x"E070",
        x"E088",
        x"E090",
        x"940E",
        x"0690",
        x"940E",
        x"0CAF",
        x"2388",
        x"F491",
        x"E184",
        x"E092",
        x"940E",
        x"1652",
        x"2D9F",
        x"2D8E",
        x"2D7D",
        x"2D6C",
        x"940E",
        x"16E2",
        x"E085",
        x"E092",
        x"940E",
        x"1652",
        x"80C9",
        x"80DA",
        x"80EB",
        x"80FC",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"16C8",
        x"06D9",
        x"06EA",
        x"06FB",
        x"F091",
        x"9180",
        x"04C3",
        x"9190",
        x"04C4",
        x"91A0",
        x"04C5",
        x"91B0",
        x"04C6",
        x"2B89",
        x"2B8A",
        x"2B8B",
        x"F081",
        x"E081",
        x"1A88",
        x"0891",
        x"08A1",
        x"08B1",
        x"F451",
        x"940E",
        x"0A4A",
        x"9080",
        x"04C3",
        x"9090",
        x"04C4",
        x"90A0",
        x"04C5",
        x"90B0",
        x"04C6",
        x"EF8F",
        x"1AC8",
        x"0AD8",
        x"0AE8",
        x"0AF8",
        x"CFAF",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"E787",
        x"E092",
        x"940E",
        x"1652",
        x"E061",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"0690",
        x"E68F",
        x"E197",
        x"9701",
        x"F7F1",
        x"C000",
        x"0000",
        x"E060",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"0690",
        x"9508",
        x"940E",
        x"0D6E",
        x"940E",
        x"0A4A",
        x"9508",
        x"E0A1",
        x"E0B0",
        x"E9E0",
        x"E0FD",
        x"940C",
        x"1AD1",
        x"8219",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17E1",
        x"E080",
        x"940E",
        x"0AAC",
        x"8189",
        x"2388",
        x"F011",
        x"940E",
        x"0D6E",
        x"EB88",
        x"E090",
        x"940E",
        x"1652",
        x"940E",
        x"0CAF",
        x"2388",
        x"F7E1",
        x"EA8B",
        x"E090",
        x"940E",
        x"1652",
        x"E081",
        x"940E",
        x"0AAC",
        x"940E",
        x"0A4A",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"0A90",
        x"FD97",
        x"C00C",
        x"2FE8",
        x"2FF9",
        x"0FEE",
        x"1FFF",
        x"51E8",
        x"4FFB",
        x"8120",
        x"8131",
        x"FF32",
        x"C002",
        x"940E",
        x"0B93",
        x"9621",
        x"E0E2",
        x"940C",
        x"1AED",
        x"E0A2",
        x"E0B0",
        x"ECEE",
        x"E0FD",
        x"940C",
        x"1ACF",
        x"9120",
        x"0299",
        x"9130",
        x"029A",
        x"3028",
        x"0531",
        x"F419",
        x"940E",
        x"0B20",
        x"C04A",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17D9",
        x"2F08",
        x"2F19",
        x"8189",
        x"819A",
        x"9601",
        x"F431",
        x"9180",
        x"0295",
        x"9190",
        x"0296",
        x"839A",
        x"8389",
        x"9180",
        x"0299",
        x"9190",
        x"029A",
        x"2F28",
        x"2F39",
        x"5F2F",
        x"4F3F",
        x"9330",
        x"029A",
        x"9320",
        x"0299",
        x"2F28",
        x"2F39",
        x"0F22",
        x"1F33",
        x"2FE2",
        x"2FF3",
        x"52E8",
        x"4FFB",
        x"8149",
        x"815A",
        x"8351",
        x"8340",
        x"2FE2",
        x"2FF3",
        x"53E9",
        x"4FFB",
        x"EF4F",
        x"EF5F",
        x"8351",
        x"8340",
        x"2FE2",
        x"2FF3",
        x"51E8",
        x"4FFB",
        x"E040",
        x"E055",
        x"8351",
        x"8340",
        x"2FE8",
        x"2FF9",
        x"54E5",
        x"4FFB",
        x"E02F",
        x"8320",
        x"940E",
        x"0B2F",
        x"2F80",
        x"2F91",
        x"940E",
        x"0D8A",
        x"9622",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"E0D0",
        x"0FCC",
        x"1FDD",
        x"2FEC",
        x"2FFD",
        x"5FEF",
        x"4FF9",
        x"95C8",
        x"2DE0",
        x"E0F0",
        x"0FEE",
        x"1FFF",
        x"5BEA",
        x"4FF9",
        x"95C8",
        x"2D00",
        x"9631",
        x"95C8",
        x"2D10",
        x"E783",
        x"E092",
        x"940E",
        x"1652",
        x"54CE",
        x"4FDF",
        x"8188",
        x"8199",
        x"940E",
        x"162D",
        x"81A8",
        x"81B9",
        x"2FEA",
        x"2FFB",
        x"9001",
        x"2000",
        x"F7E9",
        x"9731",
        x"2FCE",
        x"1BCA",
        x"30C9",
        x"F428",
        x"E280",
        x"940E",
        x"162A",
        x"5FCF",
        x"CFF9",
        x"2FE0",
        x"2FF1",
        x"95C8",
        x"2D80",
        x"2FCE",
        x"2FDF",
        x"9621",
        x"2388",
        x"F029",
        x"940E",
        x"162A",
        x"2FEC",
        x"2FFD",
        x"CFF4",
        x"E08A",
        x"940E",
        x"162A",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"2B89",
        x"F451",
        x"E78D",
        x"E094",
        x"940E",
        x"1652",
        x"9180",
        x"006D",
        x"940E",
        x"0E26",
        x"E081",
        x"9508",
        x"E080",
        x"9508",
        x"E0A5",
        x"E0B0",
        x"E8E3",
        x"E0FE",
        x"940C",
        x"1ACD",
        x"2EE6",
        x"2EF7",
        x"E041",
        x"E050",
        x"E060",
        x"E070",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"E967",
        x"E072",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6B",
        x"4F7F",
        x"940E",
        x"1801",
        x"2F08",
        x"2F19",
        x"940E",
        x"0E6F",
        x"2388",
        x"F009",
        x"C041",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"2F80",
        x"2F91",
        x"940E",
        x"1768",
        x"E683",
        x"E094",
        x"940E",
        x"1652",
        x"816D",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"0739",
        x"E08A",
        x"940E",
        x"162A",
        x"818D",
        x"940E",
        x"0757",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"940E",
        x"0768",
        x"8189",
        x"819A",
        x"81AB",
        x"81BC",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"5041",
        x"0951",
        x"0961",
        x"0971",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"1618",
        x"0619",
        x"061A",
        x"061B",
        x"F424",
        x"2DEE",
        x"2DFF",
        x"9509",
        x"CFE7",
        x"9180",
        x"0297",
        x"9190",
        x"0298",
        x"9601",
        x"9390",
        x"0298",
        x"9380",
        x"0297",
        x"9625",
        x"E0E6",
        x"940C",
        x"1AE9",
        x"EA6F",
        x"E076",
        x"940E",
        x"0E7D",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"EEEE",
        x"E0FE",
        x"940C",
        x"1ACF",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17D9",
        x"940E",
        x"0E6F",
        x"2388",
        x"F4A1",
        x"8189",
        x"819A",
        x"940E",
        x"0A90",
        x"2F08",
        x"2F19",
        x"FF97",
        x"C00F",
        x"E588",
        x"E093",
        x"940E",
        x"1652",
        x"8189",
        x"819A",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"C003",
        x"EF8F",
        x"EF9F",
        x"C002",
        x"2F80",
        x"2F91",
        x"9622",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"940E",
        x"0EE8",
        x"2F08",
        x"2F19",
        x"FD97",
        x"C021",
        x"EE8B",
        x"E090",
        x"940E",
        x"1652",
        x"2FC0",
        x"2FD1",
        x"0FCC",
        x"1FDD",
        x"2FEC",
        x"2FFD",
        x"51E8",
        x"4FFB",
        x"8180",
        x"8191",
        x"940E",
        x"0926",
        x"EE86",
        x"E090",
        x"940E",
        x"1652",
        x"52C8",
        x"4FDB",
        x"8188",
        x"8199",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"2F80",
        x"2F91",
        x"940E",
        x"0B93",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"E0A1",
        x"E0B0",
        x"E4EF",
        x"E0FF",
        x"940C",
        x"1ACF",
        x"2F08",
        x"2F19",
        x"E18F",
        x"8389",
        x"E060",
        x"E070",
        x"2F80",
        x"2F91",
        x"940E",
        x"17D9",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17E1",
        x"8189",
        x"3180",
        x"F120",
        x"ED86",
        x"E090",
        x"940E",
        x"1652",
        x"8219",
        x"8189",
        x"3180",
        x"F550",
        x"ED81",
        x"E090",
        x"940E",
        x"1652",
        x"8189",
        x"940E",
        x"166A",
        x"EC8D",
        x"E090",
        x"940E",
        x"1652",
        x"81E9",
        x"E0F0",
        x"0FEE",
        x"1FFF",
        x"5DE4",
        x"4FFE",
        x"8180",
        x"8191",
        x"940E",
        x"1652",
        x"E08A",
        x"940E",
        x"162A",
        x"8189",
        x"5F8F",
        x"8389",
        x"CFE1",
        x"2F80",
        x"2F91",
        x"940E",
        x"0EE8",
        x"FD97",
        x"C008",
        x"2FE8",
        x"2FF9",
        x"54E5",
        x"4FFB",
        x"8129",
        x"8320",
        x"940E",
        x"0B2F",
        x"9621",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"E0A5",
        x"E0B0",
        x"E9EE",
        x"E0FF",
        x"940C",
        x"1AC5",
        x"2EE6",
        x"2EF7",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"E12F",
        x"832D",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F08",
        x"2F19",
        x"940E",
        x"0E6F",
        x"2388",
        x"F009",
        x"C0D7",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"2F80",
        x"2F91",
        x"940E",
        x"17D9",
        x"2F6C",
        x"2F7D",
        x"5F6B",
        x"4F7F",
        x"940E",
        x"17E1",
        x"9180",
        x"0299",
        x"9190",
        x"029A",
        x"80AB",
        x"80BC",
        x"EDE8",
        x"E0F4",
        x"E000",
        x"E010",
        x"1708",
        x"0719",
        x"F594",
        x"9121",
        x"9131",
        x"152A",
        x"053B",
        x"F551",
        x"2FE0",
        x"2FF1",
        x"0FEE",
        x"1FFF",
        x"51E8",
        x"4FFB",
        x"8180",
        x"8191",
        x"2D2E",
        x"2D3F",
        x"2328",
        x"2339",
        x"2B23",
        x"F081",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"0926",
        x"ED85",
        x"E092",
        x"940E",
        x"1652",
        x"818B",
        x"819C",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"C099",
        x"812D",
        x"312F",
        x"F431",
        x"2FE0",
        x"2FF1",
        x"54E5",
        x"4FFB",
        x"8120",
        x"832D",
        x"2AE8",
        x"2AF9",
        x"C063",
        x"5F0F",
        x"4F1F",
        x"CFCB",
        x"1708",
        x"0719",
        x"F009",
        x"C05C",
        x"3008",
        x"0511",
        x"F419",
        x"940E",
        x"0B20",
        x"C080",
        x"818D",
        x"318F",
        x"F411",
        x"E08F",
        x"838D",
        x"2FE0",
        x"2FF1",
        x"0FEE",
        x"1FFF",
        x"2F6E",
        x"2F7F",
        x"5268",
        x"4F7B",
        x"2F2E",
        x"2F3F",
        x"5329",
        x"4F3B",
        x"2F8E",
        x"2F9F",
        x"5188",
        x"4F9B",
        x"2E68",
        x"2E79",
        x"2FA0",
        x"2FB1",
        x"54A5",
        x"4FBB",
        x"2F80",
        x"2F91",
        x"1618",
        x"0619",
        x"F04C",
        x"5F0F",
        x"4F1F",
        x"9310",
        x"029A",
        x"9300",
        x"0299",
        x"2F08",
        x"2F19",
        x"C02D",
        x"2E88",
        x"2E99",
        x"E0F1",
        x"1A8F",
        x"0891",
        x"2FE6",
        x"2FF7",
        x"90D2",
        x"90C2",
        x"2F4E",
        x"2F5F",
        x"5022",
        x"0931",
        x"E0F2",
        x"1A6F",
        x"0871",
        x"9711",
        x"14AC",
        x"04BD",
        x"F718",
        x"2FE6",
        x"2FF7",
        x"82D1",
        x"82C0",
        x"2FE2",
        x"2FF3",
        x"8180",
        x"8191",
        x"8393",
        x"8382",
        x"2DE6",
        x"2DF7",
        x"8180",
        x"8191",
        x"8393",
        x"8382",
        x"918C",
        x"9611",
        x"938C",
        x"9711",
        x"2F64",
        x"2F75",
        x"2D88",
        x"2D99",
        x"CFC7",
        x"2D6E",
        x"2D7F",
        x"818B",
        x"819C",
        x"940E",
        x"0B0A",
        x"816D",
        x"8149",
        x"815A",
        x"2F80",
        x"2F91",
        x"0F88",
        x"1F99",
        x"2FE8",
        x"2FF9",
        x"52E8",
        x"4FFB",
        x"812B",
        x"813C",
        x"2324",
        x"2335",
        x"8331",
        x"8320",
        x"2FE8",
        x"2FF9",
        x"53E9",
        x"4FFB",
        x"8351",
        x"8340",
        x"2FE8",
        x"2FF9",
        x"51E8",
        x"4FFB",
        x"82F1",
        x"82E0",
        x"2FE0",
        x"2FF1",
        x"54E5",
        x"4FFB",
        x"8360",
        x"940E",
        x"0B2F",
        x"9625",
        x"E0EE",
        x"940C",
        x"1AE1",
        x"E060",
        x"E071",
        x"940E",
        x"0F98",
        x"9508",
        x"E060",
        x"E072",
        x"940E",
        x"0F98",
        x"9508",
        x"E061",
        x"E070",
        x"940E",
        x"0F98",
        x"9508",
        x"E062",
        x"E070",
        x"940E",
        x"0F98",
        x"9508",
        x"E064",
        x"E070",
        x"940E",
        x"0F98",
        x"9508",
        x"E068",
        x"E070",
        x"940E",
        x"0F98",
        x"9508",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"921F",
        x"B7CD",
        x"B7DE",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6B",
        x"4F7F",
        x"940E",
        x"1801",
        x"940E",
        x"0E6F",
        x"2388",
        x"F5B1",
        x"EE8B",
        x"E091",
        x"940E",
        x"1652",
        x"818B",
        x"819C",
        x"940E",
        x"167A",
        x"EE86",
        x"E091",
        x"940E",
        x"1652",
        x"8189",
        x"819A",
        x"940E",
        x"167A",
        x"EE82",
        x"E091",
        x"940E",
        x"1652",
        x"818D",
        x"940E",
        x"166F",
        x"E08A",
        x"940E",
        x"162A",
        x"818D",
        x"940E",
        x"0757",
        x"818B",
        x"819C",
        x"940E",
        x"0768",
        x"80CB",
        x"80DC",
        x"2CE1",
        x"2CF1",
        x"8189",
        x"819A",
        x"E0A0",
        x"E0B0",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F044",
        x"940E",
        x"07C0",
        x"EF8F",
        x"1AC8",
        x"0AD8",
        x"0AE8",
        x"0AF8",
        x"CFEF",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"E1E5",
        x"E1F1",
        x"940C",
        x"1AD1",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17DD",
        x"940E",
        x"0E6F",
        x"2388",
        x"F479",
        x"E48C",
        x"940E",
        x"0757",
        x"8189",
        x"819A",
        x"940E",
        x"0768",
        x"E060",
        x"E070",
        x"E188",
        x"E090",
        x"940E",
        x"0690",
        x"940E",
        x"0A4A",
        x"9622",
        x"E0E2",
        x"940C",
        x"1AED",
        x"E0A3",
        x"E0B0",
        x"E3E8",
        x"E1F1",
        x"940C",
        x"1ACF",
        x"821B",
        x"821A",
        x"8219",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"1801",
        x"2F08",
        x"2F19",
        x"940E",
        x"0E6F",
        x"2388",
        x"F5A1",
        x"2F6C",
        x"2F7D",
        x"5F6E",
        x"4F7F",
        x"2F80",
        x"2F91",
        x"940E",
        x"17E1",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17E1",
        x"E080",
        x"940E",
        x"06E0",
        x"2F08",
        x"2F19",
        x"818B",
        x"940E",
        x"0757",
        x"8189",
        x"E090",
        x"2F98",
        x"2788",
        x"812A",
        x"0F82",
        x"1D91",
        x"940E",
        x"0768",
        x"E060",
        x"E070",
        x"E188",
        x"E090",
        x"940E",
        x"0690",
        x"E48C",
        x"940E",
        x"0757",
        x"2F80",
        x"2F91",
        x"940E",
        x"0768",
        x"E060",
        x"E070",
        x"E188",
        x"E090",
        x"940E",
        x"0690",
        x"940E",
        x"0A4A",
        x"9623",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17DD",
        x"940E",
        x"0E6F",
        x"2388",
        x"F5C9",
        x"818B",
        x"819C",
        x"940E",
        x"0768",
        x"808B",
        x"809C",
        x"2CA1",
        x"2CB1",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"8189",
        x"819A",
        x"E0A0",
        x"E0B0",
        x"1588",
        x"0599",
        x"05AA",
        x"05BB",
        x"F0CC",
        x"940E",
        x"06D6",
        x"E098",
        x"0CCC",
        x"1CDD",
        x"1CEE",
        x"1CFF",
        x"2F28",
        x"7021",
        x"2AC2",
        x"9586",
        x"FEE0",
        x"C004",
        x"E22D",
        x"26C2",
        x"24EE",
        x"24FF",
        x"5091",
        x"F781",
        x"EF8F",
        x"1A88",
        x"0A98",
        x"0AA8",
        x"0AB8",
        x"CFDE",
        x"ED8C",
        x"E091",
        x"940E",
        x"1652",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"E0A6",
        x"E0B0",
        x"EEEB",
        x"E1F1",
        x"940C",
        x"1ACF",
        x"2F6C",
        x"2F7D",
        x"5F6B",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17DD",
        x"940E",
        x"0E6F",
        x"2388",
        x"F4F1",
        x"E000",
        x"E010",
        x"818D",
        x"819E",
        x"812B",
        x"813C",
        x"1B28",
        x"0B39",
        x"1720",
        x"0731",
        x"F098",
        x"0F80",
        x"1F91",
        x"940E",
        x"0768",
        x"940E",
        x"06CC",
        x"940E",
        x"0757",
        x"8189",
        x"819A",
        x"0F80",
        x"1F91",
        x"940E",
        x"0768",
        x"940E",
        x"06AF",
        x"5F0F",
        x"4F1F",
        x"CFE4",
        x"9626",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"E0A6",
        x"E0B0",
        x"E2E9",
        x"E1F2",
        x"940C",
        x"1ACD",
        x"2F6C",
        x"2F7D",
        x"5F6B",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17DD",
        x"940E",
        x"0E6F",
        x"2388",
        x"F5C9",
        x"E000",
        x"E010",
        x"818D",
        x"819E",
        x"812B",
        x"813C",
        x"1B28",
        x"0B39",
        x"1720",
        x"0731",
        x"F170",
        x"0F80",
        x"1F91",
        x"940E",
        x"0768",
        x"940E",
        x"06CC",
        x"2EE8",
        x"8189",
        x"819A",
        x"0F80",
        x"1F91",
        x"940E",
        x"0768",
        x"940E",
        x"06CC",
        x"2EF8",
        x"16E8",
        x"F0C9",
        x"EC8C",
        x"E091",
        x"940E",
        x"1652",
        x"818D",
        x"819E",
        x"2D6E",
        x"0F80",
        x"1F91",
        x"940E",
        x"0739",
        x"EC88",
        x"E091",
        x"940E",
        x"1652",
        x"8189",
        x"819A",
        x"2D6F",
        x"0F80",
        x"1F91",
        x"940E",
        x"0739",
        x"E08A",
        x"940E",
        x"162A",
        x"5F0F",
        x"4F1F",
        x"CFC9",
        x"9626",
        x"E0E6",
        x"940C",
        x"1AE9",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"D000",
        x"D000",
        x"B7CD",
        x"B7DE",
        x"2F6C",
        x"2F7D",
        x"5F6D",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17DD",
        x"940E",
        x"0E6F",
        x"2388",
        x"F519",
        x"E980",
        x"E091",
        x"940E",
        x"1652",
        x"940E",
        x"1623",
        x"818B",
        x"819C",
        x"940E",
        x"0768",
        x"80CB",
        x"80DC",
        x"2CE1",
        x"2CF1",
        x"8189",
        x"819A",
        x"E0A0",
        x"E0B0",
        x"158C",
        x"059D",
        x"05AE",
        x"05BF",
        x"F054",
        x"940E",
        x"06D6",
        x"940E",
        x"160F",
        x"EF8F",
        x"1AC8",
        x"0AD8",
        x"0AE8",
        x"0AF8",
        x"CFED",
        x"940E",
        x"1623",
        x"900F",
        x"900F",
        x"900F",
        x"900F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"ECEA",
        x"E1F2",
        x"940C",
        x"1ACB",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17DD",
        x"940E",
        x"0E6F",
        x"2388",
        x"F5E1",
        x"8109",
        x"811A",
        x"940E",
        x"072C",
        x"940E",
        x"1623",
        x"940E",
        x"0757",
        x"2EC0",
        x"2ED1",
        x"EF8F",
        x"1AC8",
        x"0AD8",
        x"2F80",
        x"2F91",
        x"940E",
        x"0768",
        x"940E",
        x"06AF",
        x"EE88",
        x"2EE8",
        x"E083",
        x"2EF8",
        x"940E",
        x"1627",
        x"2388",
        x"F4F1",
        x"E68F",
        x"E197",
        x"9701",
        x"F7F1",
        x"C000",
        x"0000",
        x"E091",
        x"1AE9",
        x"08F1",
        x"F791",
        x"E889",
        x"E091",
        x"940E",
        x"1652",
        x"8189",
        x"819A",
        x"940E",
        x"167A",
        x"E884",
        x"E091",
        x"940E",
        x"1652",
        x"2F80",
        x"2F91",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"C003",
        x"2D0C",
        x"2D1D",
        x"CFC8",
        x"9622",
        x"E0E8",
        x"940C",
        x"1AE7",
        x"E0A8",
        x"E0B0",
        x"E1EA",
        x"E1F3",
        x"940C",
        x"1ACF",
        x"E94C",
        x"EF5F",
        x"EF6F",
        x"EF7F",
        x"8349",
        x"835A",
        x"836B",
        x"837C",
        x"2F6C",
        x"2F7D",
        x"5F69",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F6C",
        x"2F7D",
        x"5F6B",
        x"4F7F",
        x"940E",
        x"17DD",
        x"2F08",
        x"2F19",
        x"940E",
        x"0E6F",
        x"2388",
        x"F009",
        x"C041",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"2F80",
        x"2F91",
        x"940E",
        x"1768",
        x"8149",
        x"815A",
        x"816B",
        x"817C",
        x"812D",
        x"813E",
        x"818F",
        x"8598",
        x"394C",
        x"EFEF",
        x"075E",
        x"076E",
        x"077E",
        x"F539",
        x"E545",
        x"E050",
        x"2F62",
        x"2F73",
        x"940E",
        x"0C00",
        x"816D",
        x"817E",
        x"EA4A",
        x"E050",
        x"818F",
        x"8598",
        x"940E",
        x"0C00",
        x"816D",
        x"817E",
        x"EF4F",
        x"E050",
        x"818F",
        x"8598",
        x"940E",
        x"0C00",
        x"E000",
        x"E010",
        x"816D",
        x"817E",
        x"2F40",
        x"2F51",
        x"818F",
        x"8598",
        x"940E",
        x"0C00",
        x"5001",
        x"0911",
        x"3F08",
        x"EF8F",
        x"0718",
        x"F791",
        x"C004",
        x"2F62",
        x"2F73",
        x"940E",
        x"0C00",
        x"9628",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"E0A2",
        x"E0B0",
        x"E8E0",
        x"E1F3",
        x"940C",
        x"1ACF",
        x"839A",
        x"8389",
        x"2FE8",
        x"2FF9",
        x"8180",
        x"2388",
        x"F079",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"0634",
        x"3282",
        x"F418",
        x"940E",
        x"0E26",
        x"C024",
        x"8189",
        x"819A",
        x"940E",
        x"067E",
        x"C01F",
        x"940E",
        x"0A68",
        x"E688",
        x"E092",
        x"940E",
        x"1652",
        x"E202",
        x"E010",
        x"5F1F",
        x"EF8F",
        x"5F8F",
        x"2FE8",
        x"E0F0",
        x"0FEE",
        x"1FFF",
        x"50E0",
        x"4FFA",
        x"95C8",
        x"2DE0",
        x"23EE",
        x"F039",
        x"171E",
        x"F799",
        x"940E",
        x"0E26",
        x"5001",
        x"F769",
        x"C003",
        x"2311",
        x"F751",
        x"CFF8",
        x"9622",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2F86",
        x"940E",
        x"0757",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"0768",
        x"940E",
        x"06AF",
        x"91DF",
        x"91CF",
        x"9508",
        x"93CF",
        x"2FC8",
        x"EF6F",
        x"E483",
        x"EF9E",
        x"940E",
        x"13B9",
        x"2F6C",
        x"E48F",
        x"EF9E",
        x"940E",
        x"13B9",
        x"E060",
        x"E480",
        x"EF9E",
        x"940E",
        x"13B9",
        x"E068",
        x"E480",
        x"EF9E",
        x"940E",
        x"13B9",
        x"91CF",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FD6",
        x"2FC4",
        x"940E",
        x"13C9",
        x"2F8D",
        x"940E",
        x"13C9",
        x"2F8C",
        x"940E",
        x"13C9",
        x"91DF",
        x"91CF",
        x"9508",
        x"E0A1",
        x"E0B0",
        x"EFE6",
        x"E1F3",
        x"940C",
        x"1AC9",
        x"E027",
        x"8329",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17E1",
        x"8189",
        x"3087",
        x"F480",
        x"E090",
        x"0F88",
        x"1F99",
        x"2FE8",
        x"2FF9",
        x"5EE2",
        x"4FFE",
        x"80E0",
        x"80F1",
        x"2FE8",
        x"2FF9",
        x"5FE0",
        x"4FFE",
        x"8100",
        x"8111",
        x"C006",
        x"E000",
        x"E010",
        x"ED3E",
        x"2EE3",
        x"E034",
        x"2EF3",
        x"E06F",
        x"E482",
        x"EF9E",
        x"940E",
        x"13B9",
        x"E02F",
        x"2ED2",
        x"2D6D",
        x"E480",
        x"EF9E",
        x"940E",
        x"13B9",
        x"94DA",
        x"E027",
        x"16D2",
        x"F7B9",
        x"E98B",
        x"2EC8",
        x"E084",
        x"2ED8",
        x"EA96",
        x"2EA9",
        x"E094",
        x"2EB9",
        x"2DEC",
        x"2DFD",
        x"95C8",
        x"2D80",
        x"940E",
        x"13C9",
        x"EFFF",
        x"1ACF",
        x"0ADF",
        x"14AC",
        x"04BD",
        x"F7A1",
        x"2CD1",
        x"2D6D",
        x"E080",
        x"EF9E",
        x"940E",
        x"13B9",
        x"2DEE",
        x"2DFF",
        x"95C8",
        x"2D60",
        x"E081",
        x"EF9E",
        x"940E",
        x"13B9",
        x"94D3",
        x"EFFF",
        x"1AEF",
        x"0AFF",
        x"E120",
        x"16D2",
        x"F761",
        x"81E9",
        x"E0F0",
        x"52EA",
        x"4FFB",
        x"95C8",
        x"2D60",
        x"E280",
        x"EF9E",
        x"940E",
        x"13B9",
        x"2EE0",
        x"2EF1",
        x"E180",
        x"0EE8",
        x"1CF1",
        x"2FE0",
        x"2FF1",
        x"95C8",
        x"2D60",
        x"E281",
        x"EF9E",
        x"940E",
        x"13B9",
        x"5F0F",
        x"4F1F",
        x"150E",
        x"051F",
        x"F799",
        x"E04E",
        x"E86F",
        x"E982",
        x"940E",
        x"13E1",
        x"EFFF",
        x"E92E",
        x"E284",
        x"50F1",
        x"4020",
        x"4080",
        x"F7E1",
        x"C000",
        x"0000",
        x"E94F",
        x"E96F",
        x"E98F",
        x"940E",
        x"13E1",
        x"9621",
        x"E0EA",
        x"940C",
        x"1AE5",
        x"E0A4",
        x"E0B0",
        x"E8E9",
        x"E1F4",
        x"940C",
        x"1AD1",
        x"940E",
        x"1623",
        x"8389",
        x"940E",
        x"1623",
        x"838A",
        x"821B",
        x"2F6C",
        x"2F7D",
        x"5F6C",
        x"4F7F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"17E1",
        x"818C",
        x"9190",
        x"04D7",
        x"0F98",
        x"9390",
        x"04D7",
        x"E090",
        x"9624",
        x"E0E2",
        x"940C",
        x"1AED",
        x"E0A0",
        x"E0B0",
        x"EAEA",
        x"E1F4",
        x"940C",
        x"1AC1",
        x"940E",
        x"072C",
        x"940E",
        x"1623",
        x"2EB8",
        x"2CC1",
        x"2CD1",
        x"24EE",
        x"94EA",
        x"2CFE",
        x"E000",
        x"E010",
        x"E0C0",
        x"E0D0",
        x"2C81",
        x"2C91",
        x"E583",
        x"16B8",
        x"F409",
        x"C040",
        x"24AA",
        x"94AA",
        x"2CBA",
        x"940E",
        x"1627",
        x"2388",
        x"F009",
        x"C08E",
        x"E081",
        x"1AA8",
        x"08B1",
        x"F7B9",
        x"E78A",
        x"E091",
        x"940E",
        x"1652",
        x"2D88",
        x"2D99",
        x"940E",
        x"16C0",
        x"E68A",
        x"E091",
        x"940E",
        x"1652",
        x"2F8C",
        x"2F9D",
        x"940E",
        x"16C0",
        x"E58C",
        x"E091",
        x"940E",
        x"1652",
        x"E48D",
        x"E091",
        x"940E",
        x"1652",
        x"2F80",
        x"2F91",
        x"940E",
        x"167A",
        x"E480",
        x"E091",
        x"940E",
        x"1652",
        x"2D8E",
        x"2D9F",
        x"940E",
        x"167A",
        x"E38A",
        x"E091",
        x"940E",
        x"1652",
        x"2D8C",
        x"2D9D",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"B7CD",
        x"B7DE",
        x"E1E2",
        x"940C",
        x"1ADD",
        x"940E",
        x"1623",
        x"2EB8",
        x"E381",
        x"16B8",
        x"F059",
        x"E28F",
        x"E091",
        x"940E",
        x"1652",
        x"2D8B",
        x"940E",
        x"162A",
        x"E08A",
        x"940E",
        x"162A",
        x"CFAB",
        x"E081",
        x"9380",
        x"04D7",
        x"940E",
        x"1483",
        x"2E38",
        x"EF8D",
        x"2E28",
        x"0C23",
        x"940E",
        x"1483",
        x"2EB8",
        x"940E",
        x"1483",
        x"2C7B",
        x"2C61",
        x"2C46",
        x"2C57",
        x"0E48",
        x"1E59",
        x"E083",
        x"1638",
        x"F0E9",
        x"940E",
        x"1483",
        x"144E",
        x"045F",
        x"F410",
        x"2CE4",
        x"2CF5",
        x"14C4",
        x"04D5",
        x"F410",
        x"2CC4",
        x"2CD5",
        x"940E",
        x"0757",
        x"2CA4",
        x"2CB5",
        x"EF8F",
        x"1AA8",
        x"0AB8",
        x"2D84",
        x"2D95",
        x"940E",
        x"0768",
        x"940E",
        x"07C0",
        x"943A",
        x"2C4A",
        x"2C5B",
        x"CFE0",
        x"0D02",
        x"1D11",
        x"940E",
        x"1483",
        x"940E",
        x"1623",
        x"2EB8",
        x"9180",
        x"04D7",
        x"2388",
        x"F011",
        x"9621",
        x"CF6A",
        x"EF8F",
        x"1A88",
        x"0A98",
        x"CF66",
        x"940E",
        x"1623",
        x"2EB8",
        x"CF62",
        x"93CF",
        x"2FC6",
        x"940E",
        x"162D",
        x"23CC",
        x"F019",
        x"E283",
        x"E091",
        x"C002",
        x"E189",
        x"E091",
        x"940E",
        x"1652",
        x"91CF",
        x"9508",
        x"E0A1",
        x"E0B0",
        x"E6ED",
        x"E1F5",
        x"940C",
        x"1AD1",
        x"EF2F",
        x"8329",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"17E1",
        x"8189",
        x"3084",
        x"F440",
        x"B398",
        x"739F",
        x"9582",
        x"0F88",
        x"0F88",
        x"7C80",
        x"2B89",
        x"BB88",
        x"B368",
        x"7860",
        x"E689",
        x"E091",
        x"940E",
        x"1558",
        x"B368",
        x"7460",
        x"E68D",
        x"E091",
        x"940E",
        x"1558",
        x"9621",
        x"E0E2",
        x"940C",
        x"1AED",
        x"BA1A",
        x"EF8F",
        x"BB87",
        x"E38F",
        x"BB81",
        x"B812",
        x"BA18",
        x"E060",
        x"EC72",
        x"E081",
        x"E090",
        x"940E",
        x"1643",
        x"940E",
        x"0A68",
        x"940E",
        x"0B2F",
        x"E060",
        x"E070",
        x"E086",
        x"E090",
        x"940E",
        x"0690",
        x"E060",
        x"E070",
        x"E08A",
        x"E090",
        x"940E",
        x"0690",
        x"E081",
        x"940E",
        x"0AAC",
        x"E061",
        x"E070",
        x"E080",
        x"E090",
        x"940E",
        x"0AB7",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"EBED",
        x"E1F5",
        x"940C",
        x"1AD1",
        x"839A",
        x"8389",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"0634",
        x"2FE8",
        x"8189",
        x"819A",
        x"2FA8",
        x"2FB9",
        x"912C",
        x"332F",
        x"F421",
        x"2F8E",
        x"940E",
        x"0E26",
        x"C010",
        x"32E2",
        x"F460",
        x"93E0",
        x"006D",
        x"E0F0",
        x"0FEE",
        x"1FFF",
        x"59E2",
        x"4FFF",
        x"9001",
        x"81F0",
        x"2DE0",
        x"9509",
        x"C002",
        x"940E",
        x"067E",
        x"9622",
        x"E0E2",
        x"940C",
        x"1AED",
        x"9180",
        x"0294",
        x"2388",
        x"F0A9",
        x"EA86",
        x"E090",
        x"940E",
        x"1652",
        x"9180",
        x"0294",
        x"FF80",
        x"C003",
        x"E988",
        x"E090",
        x"C004",
        x"FF81",
        x"C004",
        x"E889",
        x"E090",
        x"940E",
        x"1652",
        x"E883",
        x"E090",
        x"940E",
        x"1652",
        x"9210",
        x"0294",
        x"9508",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"E188",
        x"B98A",
        x"E660",
        x"EE73",
        x"E186",
        x"E090",
        x"940E",
        x"1A8F",
        x"5021",
        x"B929",
        x"9508",
        x"9B5D",
        x"CFFE",
        x"B98C",
        x"9508",
        x"308D",
        x"F011",
        x"308A",
        x"F421",
        x"E08D",
        x"940E",
        x"160F",
        x"E08A",
        x"940E",
        x"160F",
        x"9508",
        x"940E",
        x"1613",
        x"E080",
        x"E090",
        x"9508",
        x"9B5F",
        x"CFFE",
        x"B18C",
        x"9508",
        x"B18B",
        x"7880",
        x"9508",
        x"940E",
        x"1613",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"9189",
        x"2388",
        x"F019",
        x"940E",
        x"1613",
        x"CFFA",
        x"91DF",
        x"91CF",
        x"9508",
        x"E887",
        x"E092",
        x"940E",
        x"162D",
        x"E88C",
        x"E092",
        x"940E",
        x"162D",
        x"9508",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F429",
        x"E188",
        x"B98A",
        x"E98B",
        x"B989",
        x"C002",
        x"940E",
        x"1600",
        x"940E",
        x"163A",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2FEC",
        x"2FFD",
        x"95C8",
        x"2D80",
        x"2388",
        x"F021",
        x"9621",
        x"940E",
        x"1613",
        x"CFF6",
        x"91DF",
        x"91CF",
        x"9508",
        x"708F",
        x"308A",
        x"F410",
        x"5D80",
        x"9508",
        x"5C89",
        x"9508",
        x"940E",
        x"1663",
        x"940E",
        x"1613",
        x"9508",
        x"93CF",
        x"2FC8",
        x"9582",
        x"708F",
        x"940E",
        x"166A",
        x"2F8C",
        x"940E",
        x"166A",
        x"91CF",
        x"9508",
        x"93CF",
        x"2FC8",
        x"2F89",
        x"940E",
        x"166F",
        x"2F8C",
        x"940E",
        x"166F",
        x"91CF",
        x"9508",
        x"2F28",
        x"2F39",
        x"2FE8",
        x"2FF9",
        x"2F94",
        x"5091",
        x"F010",
        x"9361",
        x"CFFC",
        x"2F82",
        x"2F93",
        x"0F84",
        x"1D91",
        x"9508",
        x"93CF",
        x"93DF",
        x"2FD8",
        x"2FC9",
        x"2F86",
        x"940E",
        x"1663",
        x"2FED",
        x"2FFC",
        x"9381",
        x"2F8E",
        x"2F9F",
        x"91DF",
        x"91CF",
        x"9508",
        x"93CF",
        x"2FC6",
        x"9562",
        x"706F",
        x"940E",
        x"1692",
        x"2F6C",
        x"940E",
        x"1692",
        x"91CF",
        x"9508",
        x"93CF",
        x"2FC6",
        x"2F67",
        x"940E",
        x"16A1",
        x"2F6C",
        x"940E",
        x"16A1",
        x"91CF",
        x"9508",
        x"2F28",
        x"2F39",
        x"2F86",
        x"2F97",
        x"E04A",
        x"2F62",
        x"2F73",
        x"940E",
        x"1B84",
        x"9508",
        x"E1A0",
        x"E0B0",
        x"ECE6",
        x"E1F6",
        x"940C",
        x"1AD1",
        x"2F68",
        x"2F79",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"16B6",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"162D",
        x"9660",
        x"E0E2",
        x"940C",
        x"1AED",
        x"2FE8",
        x"2FF9",
        x"2F97",
        x"2F86",
        x"2F75",
        x"2F64",
        x"E02A",
        x"2F4E",
        x"2F5F",
        x"940E",
        x"1B8F",
        x"9508",
        x"E1A0",
        x"E0B0",
        x"EEE8",
        x"E1F6",
        x"940C",
        x"1AD1",
        x"2F46",
        x"2F57",
        x"2F68",
        x"2F79",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"16D6",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"162D",
        x"9660",
        x"E0E2",
        x"940C",
        x"1AED",
        x"2FE6",
        x"2FF7",
        x"9121",
        x"2F6E",
        x"2F7F",
        x"2322",
        x"F031",
        x"2FE8",
        x"2FF9",
        x"9321",
        x"2F8E",
        x"2F9F",
        x"CFF3",
        x"9508",
        x"E99F",
        x"0F98",
        x"3096",
        x"F410",
        x"5287",
        x"C005",
        x"EB9F",
        x"0F98",
        x"3096",
        x"F408",
        x"5087",
        x"ED90",
        x"0F98",
        x"3190",
        x"F410",
        x"708F",
        x"9508",
        x"EF8F",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"E2E1",
        x"E1F7",
        x"940C",
        x"1AC8",
        x"9700",
        x"F199",
        x"2FC8",
        x"2FD9",
        x"2ECC",
        x"2EDD",
        x"2F2C",
        x"2F3D",
        x"5F2F",
        x"4F3F",
        x"8188",
        x"3280",
        x"F419",
        x"2FC2",
        x"2FD3",
        x"CFF4",
        x"2E94",
        x"2EA6",
        x"2EB7",
        x"2CE1",
        x"2CF1",
        x"2F0C",
        x"2F1D",
        x"9621",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"940E",
        x"1708",
        x"FD87",
        x"C011",
        x"E094",
        x"0CEE",
        x"1CFF",
        x"959A",
        x"F7E1",
        x"0EE8",
        x"1CF1",
        x"FD87",
        x"94FA",
        x"14A1",
        x"04B1",
        x"F351",
        x"2DEA",
        x"2DFB",
        x"82F1",
        x"82E0",
        x"CFE5",
        x"2099",
        x"F031",
        x"16C0",
        x"06D1",
        x"F419",
        x"E080",
        x"E090",
        x"C002",
        x"2F80",
        x"2F91",
        x"B7CD",
        x"B7DE",
        x"E0EB",
        x"940C",
        x"1AE4",
        x"ED90",
        x"0F98",
        x"309A",
        x"F410",
        x"708F",
        x"9508",
        x"EF8F",
        x"9508",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"2EA6",
        x"2EB7",
        x"2B89",
        x"F409",
        x"C049",
        x"2FEC",
        x"2FFD",
        x"8188",
        x"9621",
        x"3280",
        x"F3D1",
        x"328D",
        x"F421",
        x"2FEC",
        x"2FFD",
        x"EF8F",
        x"C001",
        x"E081",
        x"2F0E",
        x"2F1F",
        x"2CC1",
        x"2CD1",
        x"2CE1",
        x"2CF1",
        x"2E48",
        x"0F88",
        x"0855",
        x"0866",
        x"0877",
        x"2FC0",
        x"2FD1",
        x"5F0F",
        x"4F1F",
        x"8188",
        x"940E",
        x"1708",
        x"2E98",
        x"FD87",
        x"C027",
        x"E02A",
        x"E030",
        x"E040",
        x"E050",
        x"2D9F",
        x"2D8E",
        x"2D7D",
        x"2D6C",
        x"940E",
        x"1A74",
        x"2CC9",
        x"0C99",
        x"08DD",
        x"08EE",
        x"08FF",
        x"0EC6",
        x"1ED7",
        x"1EE8",
        x"1EF9",
        x"14A1",
        x"04B1",
        x"F301",
        x"2D5F",
        x"2D4E",
        x"2D3D",
        x"2D2C",
        x"2D97",
        x"2D86",
        x"2D75",
        x"2D64",
        x"940E",
        x"1A74",
        x"2DEA",
        x"2DFB",
        x"8360",
        x"8371",
        x"8382",
        x"8393",
        x"CFCF",
        x"2F8C",
        x"2F9D",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"907F",
        x"906F",
        x"905F",
        x"904F",
        x"9508",
        x"E040",
        x"940E",
        x"171B",
        x"9508",
        x"E041",
        x"940E",
        x"171B",
        x"9508",
        x"E0A2",
        x"E0B0",
        x"EEE7",
        x"E1F7",
        x"940C",
        x"1ACF",
        x"2F06",
        x"2F17",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"E040",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"171B",
        x"8129",
        x"813A",
        x"3F2F",
        x"EF4F",
        x"0734",
        x"F019",
        x"2FE0",
        x"2FF1",
        x"8320",
        x"9622",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"E0A2",
        x"E0B0",
        x"E0E7",
        x"E1F8",
        x"940C",
        x"1ACF",
        x"2F06",
        x"2F17",
        x"EF2F",
        x"EF3F",
        x"833A",
        x"8329",
        x"E041",
        x"2F6C",
        x"2F7D",
        x"5F6F",
        x"4F7F",
        x"940E",
        x"171B",
        x"8129",
        x"813A",
        x"3F2F",
        x"EF4F",
        x"0734",
        x"F019",
        x"2FE0",
        x"2FF1",
        x"8320",
        x"9622",
        x"E0E4",
        x"940C",
        x"1AEB",
        x"92AF",
        x"92BF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"97A8",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2EE8",
        x"2EF9",
        x"940E",
        x"06D6",
        x"2F18",
        x"2EA8",
        x"2CB1",
        x"2DEA",
        x"2DFB",
        x"55E1",
        x"4FF8",
        x"95C8",
        x"2D00",
        x"E248",
        x"E260",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"1684",
        x"E38A",
        x"838E",
        x"8B89",
        x"2D6E",
        x"2D7F",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"16AC",
        x"2F61",
        x"2F8C",
        x"2F9D",
        x"9608",
        x"940E",
        x"16A1",
        x"3003",
        x"F428",
        x"EF8F",
        x"1AE8",
        x"0AF8",
        x"E010",
        x"C00E",
        x"940E",
        x"06D6",
        x"2F18",
        x"2F68",
        x"2F8C",
        x"2F9D",
        x"960B",
        x"940E",
        x"16A1",
        x"300C",
        x"F428",
        x"E0A2",
        x"0EEA",
        x"1CF1",
        x"2CD1",
        x"C00C",
        x"940E",
        x"06D6",
        x"2ED8",
        x"2F68",
        x"2F8C",
        x"2F9D",
        x"960E",
        x"940E",
        x"16A1",
        x"E0B3",
        x"0EEB",
        x"1CF1",
        x"2DEA",
        x"2DFB",
        x"55E1",
        x"4FF7",
        x"95C8",
        x"2D80",
        x"E090",
        x"E063",
        x"E070",
        x"940E",
        x"1A63",
        x"2FAC",
        x"2FBD",
        x"9653",
        x"E020",
        x"E030",
        x"2FE8",
        x"2FF9",
        x"0FE2",
        x"1FF3",
        x"55E1",
        x"4FF6",
        x"95C8",
        x"2DE0",
        x"93ED",
        x"5F2F",
        x"4F3F",
        x"3023",
        x"0531",
        x"F791",
        x"2F40",
        x"E050",
        x"2FE4",
        x"2FF5",
        x"9731",
        x"31E0",
        x"05F1",
        x"F008",
        x"C0D0",
        x"5DE0",
        x"4FFF",
        x"940C",
        x"1AB6",
        x"E481",
        x"8B8F",
        x"2FEC",
        x"2FFD",
        x"9678",
        x"C0C9",
        x"E284",
        x"8B8F",
        x"2D6E",
        x"2D7F",
        x"0F61",
        x"1D71",
        x"FD17",
        x"957A",
        x"2F8C",
        x"2F9D",
        x"9648",
        x"940E",
        x"16AC",
        x"C011",
        x"E283",
        x"8B8F",
        x"2F8C",
        x"2F9D",
        x"9648",
        x"C003",
        x"2F8C",
        x"2F9D",
        x"9647",
        x"E224",
        x"2FE8",
        x"2FF9",
        x"8320",
        x"2F61",
        x"9601",
        x"940E",
        x"16A1",
        x"2FE8",
        x"2FF9",
        x"C0A7",
        x"E284",
        x"8B8F",
        x"2F61",
        x"2F8C",
        x"2F9D",
        x"9648",
        x"940E",
        x"16A1",
        x"E22C",
        x"2FA8",
        x"2FB9",
        x"932C",
        x"2FE8",
        x"2FF9",
        x"9632",
        x"E528",
        x"C05F",
        x"E284",
        x"8B8F",
        x"2F61",
        x"2F8C",
        x"2F9D",
        x"9648",
        x"C04E",
        x"E288",
        x"8B8F",
        x"E284",
        x"8F88",
        x"2F61",
        x"2F8C",
        x"2F9D",
        x"9649",
        x"C05D",
        x"E288",
        x"8B8F",
        x"E284",
        x"8F88",
        x"2F61",
        x"2F8C",
        x"2F9D",
        x"9649",
        x"C069",
        x"E288",
        x"8B8F",
        x"E284",
        x"8F88",
        x"2F61",
        x"2F8C",
        x"2F9D",
        x"9649",
        x"940E",
        x"16A1",
        x"2FA8",
        x"2FB9",
        x"E289",
        x"938C",
        x"E28C",
        x"9611",
        x"938C",
        x"9711",
        x"2FEA",
        x"2FFB",
        x"9633",
        x"E589",
        x"C060",
        x"E284",
        x"8B8F",
        x"2D6D",
        x"2F8C",
        x"2F9D",
        x"9648",
        x"940E",
        x"16A1",
        x"2F61",
        x"CFB0",
        x"E284",
        x"8B8F",
        x"2D6D",
        x"2F8C",
        x"2F9D",
        x"9648",
        x"940E",
        x"16A1",
        x"2F61",
        x"940E",
        x"16A1",
        x"E22C",
        x"2FE8",
        x"2FF9",
        x"8320",
        x"9632",
        x"E528",
        x"C011",
        x"E284",
        x"8B8F",
        x"2D6D",
        x"2F8C",
        x"2F9D",
        x"9648",
        x"940E",
        x"16A1",
        x"2F61",
        x"940E",
        x"16A1",
        x"E22C",
        x"2FE8",
        x"2FF9",
        x"8320",
        x"9632",
        x"E529",
        x"2FA8",
        x"2FB9",
        x"9611",
        x"932C",
        x"C034",
        x"E288",
        x"8B8F",
        x"E284",
        x"8F88",
        x"2D6D",
        x"2F8C",
        x"2F9D",
        x"9649",
        x"940E",
        x"16A1",
        x"2F61",
        x"940E",
        x"16A1",
        x"2FE8",
        x"2FF9",
        x"9631",
        x"E229",
        x"2FA8",
        x"2FB9",
        x"932C",
        x"C01F",
        x"E288",
        x"8B8F",
        x"E284",
        x"8F88",
        x"2D6D",
        x"2F8C",
        x"2F9D",
        x"9649",
        x"940E",
        x"16A1",
        x"2F61",
        x"940E",
        x"16A1",
        x"2FA8",
        x"2FB9",
        x"E28C",
        x"938C",
        x"E588",
        x"9611",
        x"938C",
        x"9711",
        x"2FEA",
        x"2FFB",
        x"9633",
        x"E289",
        x"9612",
        x"938C",
        x"C003",
        x"2FEC",
        x"2FFD",
        x"9677",
        x"E08A",
        x"8380",
        x"8211",
        x"2F8C",
        x"2F9D",
        x"9601",
        x"940E",
        x"162D",
        x"2D8E",
        x"2D9F",
        x"96A8",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90BF",
        x"90AF",
        x"9508",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"E283",
        x"940E",
        x"06C1",
        x"2FC8",
        x"E0D0",
        x"E988",
        x"E09A",
        x"940E",
        x"1652",
        x"E280",
        x"940E",
        x"06C1",
        x"940E",
        x"166F",
        x"E984",
        x"E09A",
        x"940E",
        x"1652",
        x"E281",
        x"940E",
        x"06C1",
        x"940E",
        x"166F",
        x"E980",
        x"E09A",
        x"940E",
        x"1652",
        x"E282",
        x"940E",
        x"06C1",
        x"940E",
        x"166F",
        x"E889",
        x"E09A",
        x"940E",
        x"1652",
        x"E284",
        x"940E",
        x"06C1",
        x"940E",
        x"166F",
        x"E884",
        x"E09A",
        x"940E",
        x"1652",
        x"E286",
        x"940E",
        x"06E0",
        x"940E",
        x"167A",
        x"E08A",
        x"940E",
        x"162A",
        x"E789",
        x"E09A",
        x"940E",
        x"1652",
        x"E004",
        x"E011",
        x"FFC7",
        x"C004",
        x"2FE0",
        x"2FF1",
        x"8180",
        x"C001",
        x"E28D",
        x"940E",
        x"162A",
        x"0FCC",
        x"1FDD",
        x"5F0F",
        x"4F1F",
        x"E0F1",
        x"300C",
        x"071F",
        x"F779",
        x"E08A",
        x"940E",
        x"162A",
        x"91DF",
        x"91CF",
        x"911F",
        x"910F",
        x"9508",
        x"940E",
        x"1590",
        x"940E",
        x"15E4",
        x"E080",
        x"E090",
        x"940E",
        x"0D8A",
        x"E0D0",
        x"EFCF",
        x"940E",
        x"15E4",
        x"2F6D",
        x"E98B",
        x"E092",
        x"940E",
        x"05B9",
        x"2FD8",
        x"2388",
        x"F1A9",
        x"FFC7",
        x"C007",
        x"FF87",
        x"C064",
        x"91C0",
        x"0060",
        x"FFC7",
        x"C01D",
        x"C05F",
        x"2F8C",
        x"0F8D",
        x"708F",
        x"9190",
        x"0060",
        x"FFD7",
        x"C011",
        x"1789",
        x"F099",
        x"2FE8",
        x"2E08",
        x"0C00",
        x"0BFF",
        x"E055",
        x"0FEE",
        x"1FFF",
        x"955A",
        x"F7E1",
        x"54E5",
        x"4FFD",
        x"8190",
        x"2399",
        x"F029",
        x"C003",
        x"17C9",
        x"F409",
        x"C043",
        x"2FC8",
        x"2F6C",
        x"2E0C",
        x"0C00",
        x"0B77",
        x"E045",
        x"0F66",
        x"1F77",
        x"954A",
        x"F7E1",
        x"5465",
        x"4F7D",
        x"E98B",
        x"E092",
        x"940E",
        x"1B6B",
        x"CFC1",
        x"9180",
        x"029B",
        x"2388",
        x"F409",
        x"CFBB",
        x"91C0",
        x"0060",
        x"FDC7",
        x"C011",
        x"2F8C",
        x"2E0C",
        x"0C00",
        x"0B99",
        x"E035",
        x"0F88",
        x"1F99",
        x"953A",
        x"F7E1",
        x"E96B",
        x"E072",
        x"5485",
        x"4F9D",
        x"940E",
        x"1B60",
        x"2B89",
        x"F099",
        x"E081",
        x"0F8C",
        x"708F",
        x"9380",
        x"0060",
        x"2E08",
        x"0C00",
        x"0B99",
        x"E025",
        x"0F88",
        x"1F99",
        x"952A",
        x"F7E1",
        x"E96B",
        x"E072",
        x"5485",
        x"4F9D",
        x"940E",
        x"1B6B",
        x"E98B",
        x"E092",
        x"940E",
        x"15B7",
        x"CF8E",
        x"EFCF",
        x"E0D0",
        x"CF8C",
        x"2400",
        x"2755",
        x"C004",
        x"0E08",
        x"1F59",
        x"0F88",
        x"1F99",
        x"9700",
        x"F029",
        x"9576",
        x"9567",
        x"F3B8",
        x"0571",
        x"F7B9",
        x"2D80",
        x"2F95",
        x"9508",
        x"27EE",
        x"27FF",
        x"27AA",
        x"27BB",
        x"C008",
        x"0FA2",
        x"1FB3",
        x"1FE4",
        x"1FF5",
        x"0F22",
        x"1F33",
        x"1F44",
        x"1F55",
        x"9596",
        x"9587",
        x"9577",
        x"9567",
        x"F398",
        x"4070",
        x"F7A9",
        x"9700",
        x"F799",
        x"2F6A",
        x"2F7B",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"E2A1",
        x"2E1A",
        x"1BAA",
        x"1BBB",
        x"2FEA",
        x"2FFB",
        x"C00D",
        x"1FAA",
        x"1FBB",
        x"1FEE",
        x"1FFF",
        x"17A2",
        x"07B3",
        x"07E4",
        x"07F5",
        x"F020",
        x"1BA2",
        x"0BB3",
        x"0BE4",
        x"0BF5",
        x"1F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"941A",
        x"F769",
        x"9560",
        x"9570",
        x"9580",
        x"9590",
        x"2F26",
        x"2F37",
        x"2F48",
        x"2F59",
        x"2F6A",
        x"2F7B",
        x"2F8E",
        x"2F9F",
        x"9508",
        x"0FEE",
        x"1FFF",
        x"2400",
        x"1C00",
        x"BE0B",
        x"95D8",
        x"920F",
        x"9631",
        x"95D8",
        x"920F",
        x"9508",
        x"922F",
        x"923F",
        x"924F",
        x"925F",
        x"926F",
        x"927F",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"930F",
        x"931F",
        x"93CF",
        x"93DF",
        x"B7CD",
        x"B7DE",
        x"1BCA",
        x"0BDB",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"9409",
        x"882A",
        x"8839",
        x"8848",
        x"845F",
        x"846E",
        x"847D",
        x"848C",
        x"849B",
        x"84AA",
        x"84B9",
        x"84C8",
        x"80DF",
        x"80EE",
        x"80FD",
        x"810C",
        x"811B",
        x"81AA",
        x"81B9",
        x"0FCE",
        x"1DD1",
        x"B60F",
        x"94F8",
        x"BFDE",
        x"BE0F",
        x"BFCD",
        x"2FCA",
        x"2FDB",
        x"9508",
        x"928F",
        x"929F",
        x"92AF",
        x"92BF",
        x"92CF",
        x"92DF",
        x"92EF",
        x"92FF",
        x"93CF",
        x"93DF",
        x"2FC8",
        x"2FD9",
        x"8168",
        x"8179",
        x"818A",
        x"819B",
        x"1561",
        x"0571",
        x"0581",
        x"0591",
        x"F421",
        x"E264",
        x"ED79",
        x"E58B",
        x"E097",
        x"E12D",
        x"EF33",
        x"E041",
        x"E050",
        x"940E",
        x"1BF0",
        x"2E82",
        x"2E93",
        x"2EA4",
        x"2EB5",
        x"EA27",
        x"E431",
        x"E040",
        x"E050",
        x"940E",
        x"1A74",
        x"2EC6",
        x"2ED7",
        x"2EE8",
        x"2EF9",
        x"EE2C",
        x"EF34",
        x"EF4F",
        x"EF5F",
        x"2D9B",
        x"2D8A",
        x"2D79",
        x"2D68",
        x"940E",
        x"1A74",
        x"2FB9",
        x"2FA8",
        x"2F97",
        x"2F86",
        x"0D8C",
        x"1D9D",
        x"1DAE",
        x"1DBF",
        x"FFB7",
        x"C003",
        x"9701",
        x"09A1",
        x"48B0",
        x"8388",
        x"8399",
        x"83AA",
        x"83BB",
        x"779F",
        x"91DF",
        x"91CF",
        x"90FF",
        x"90EF",
        x"90DF",
        x"90CF",
        x"90BF",
        x"90AF",
        x"909F",
        x"908F",
        x"9508",
        x"940E",
        x"1AF9",
        x"9508",
        x"E08C",
        x"E091",
        x"940E",
        x"1AF9",
        x"9508",
        x"E0A0",
        x"E0B0",
        x"9380",
        x"010C",
        x"9390",
        x"010D",
        x"93A0",
        x"010E",
        x"93B0",
        x"010F",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"918D",
        x"9001",
        x"1980",
        x"1001",
        x"F3D9",
        x"0B99",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"9001",
        x"920D",
        x"2000",
        x"F7E1",
        x"9508",
        x"2FE6",
        x"2FF7",
        x"2FA8",
        x"2FB9",
        x"5041",
        x"4050",
        x"F030",
        x"918D",
        x"9001",
        x"1980",
        x"F419",
        x"2000",
        x"F7B9",
        x"1B88",
        x"0B99",
        x"9508",
        x"27BB",
        x"304A",
        x"F431",
        x"2399",
        x"F422",
        x"E2BD",
        x"9590",
        x"9581",
        x"4F9F",
        x"940C",
        x"1BC3",
        x"27BB",
        x"302A",
        x"F451",
        x"2399",
        x"F442",
        x"E2BD",
        x"9590",
        x"9580",
        x"9570",
        x"9561",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"940C",
        x"1B9F",
        x"27BB",
        x"2FE4",
        x"2FF5",
        x"2FA6",
        x"1762",
        x"0571",
        x"0581",
        x"0591",
        x"0B33",
        x"FB30",
        x"F066",
        x"27AA",
        x"0F66",
        x"1F77",
        x"1F88",
        x"1F99",
        x"1FAA",
        x"17A2",
        x"F010",
        x"1BA2",
        x"9563",
        x"5038",
        x"F7A9",
        x"5DA0",
        x"33AA",
        x"F008",
        x"5DA9",
        x"93A1",
        x"F736",
        x"11B1",
        x"93B1",
        x"8210",
        x"2F84",
        x"2F95",
        x"940C",
        x"1BDE",
        x"27BB",
        x"2FE6",
        x"2FF7",
        x"2755",
        x"27AA",
        x"0F88",
        x"1F99",
        x"1FAA",
        x"17A4",
        x"F010",
        x"1BA4",
        x"9583",
        x"5150",
        x"F7B9",
        x"5DA0",
        x"33AA",
        x"F008",
        x"5DA9",
        x"93A1",
        x"9700",
        x"F779",
        x"11B1",
        x"93B1",
        x"9211",
        x"2F86",
        x"2F97",
        x"940C",
        x"1BDE",
        x"2FA8",
        x"2FB9",
        x"2FE8",
        x"2FF9",
        x"2F67",
        x"9171",
        x"2377",
        x"F7E1",
        x"9732",
        x"C004",
        x"917C",
        x"936D",
        x"8370",
        x"9162",
        x"17AE",
        x"07BF",
        x"F3C8",
        x"9508",
        x"2E05",
        x"FB97",
        x"F41E",
        x"9400",
        x"940E",
        x"1C07",
        x"FD57",
        x"D007",
        x"940E",
        x"1A8F",
        x"FC07",
        x"D003",
        x"F44E",
        x"940C",
        x"1C07",
        x"9550",
        x"9540",
        x"9530",
        x"9521",
        x"4F3F",
        x"4F4F",
        x"4F5F",
        x"9508",
        x"9590",
        x"9580",
        x"9570",
        x"9561",
        x"4F7F",
        x"4F8F",
        x"4F9F",
        x"9508",
        x"94F8",
        x"CFFF",
        x"71FF",
        x"7701",
        x"8401",
        x"9901",
        x"A901",
        x"C101",
        x"FF01",
        x"057B",
        x"137A",
        x"0D8A",
        x"0DC8",
        x"0CC9",
        x"198D",
        x"077E",
        x"06B6",
        x"10AC",
        x"117F",
        x"11E5",
        x"1223",
        x"085F",
        x"08D6",
        x"0EE3",
        x"110F",
        x"1132",
        x"13F0",
        x"1314",
        x"12C4",
        x"127C",
        x"14A4",
        x"1567",
        x"0D85",
        x"0AE8",
        x"0964",
        x"108E",
        x"1093",
        x"1098",
        x"109D",
        x"10A2",
        x"10A7",
        x"0F19",
        x"0F49",
        x"01C8",
        x"01D0",
        x"01D5",
        x"01DE",
        x"01E3",
        x"01E8",
        x"01ED",
        x"01F1",
        x"01F7",
        x"01FC",
        x"0200",
        x"0205",
        x"020D",
        x"0181",
        x"0211",
        x"0214",
        x"0217",
        x"021C",
        x"0221",
        x"0226",
        x"022B",
        x"0230",
        x"0235",
        x"023D",
        x"0243",
        x"0249",
        x"024F",
        x"0256",
        x"025D",
        x"0264",
        x"026B",
        x"0272",
        x"0279",
        x"027F",
        x"0000",
        x"0200",
        x"0000",
        x"0000",
        x"161E",
        x"0000",
        x"0000",
        x"564E",
        x"422D",
        x"4944",
        x"435A",
        x"0001",
        x"0000",
        x"04C6",
        x"04B6",
        x"04A6",
        x"04C6",
        x"04C6",
        x"04B6",
        x"04C6",
        x"051E",
        x"051E",
        x"051E",
        x"050E",
        x"04FE",
        x"04FE",
        x"04EE",
        x"057A",
        x"056E",
        x"056F",
        x"0576",
        x"0563",
        x"055F",
        x"0555",
        x"054A",
        x"0564",
        x"053F",
        x"0560",
        x"054B",
        x"056B",
        x"0535",
        x"0536",
        x"052E",
        x"05F3",
        x"05E6",
        x"05D9",
        x"05CC",
        x"05C0",
        x"05B4",
        x"05A8",
        x"059C",
        x"0593",
        x"058A",
        x"0580",
        x"3A20",
        x"0020",
        x"2820",
        x"4E00",
        x"494D",
        x"4900",
        x"5152",
        x"4600",
        x"7869",
        x"6465",
        x"4300",
        x"6568",
        x"6B63",
        x"7265",
        x"6F62",
        x"7261",
        x"0064",
        x"6E49",
        x"6576",
        x"7372",
        x"2065",
        x"6863",
        x"6365",
        x"656B",
        x"6272",
        x"616F",
        x"6472",
        x"4100",
        x"6464",
        x"6572",
        x"7373",
        x"7020",
        x"7461",
        x"6574",
        x"6E72",
        x"4900",
        x"766E",
        x"7265",
        x"6573",
        x"6120",
        x"6464",
        x"6572",
        x"7373",
        x"7020",
        x"7461",
        x"6574",
        x"6E72",
        x"5200",
        x"6E61",
        x"6F64",
        x"006D",
        x"6968",
        x"7473",
        x"726F",
        x"0079",
        x"6568",
        x"706C",
        x"6300",
        x"6E6F",
        x"6974",
        x"756E",
        x"0065",
        x"656E",
        x"7478",
        x"7300",
        x"6574",
        x"0070",
        x"6572",
        x"7367",
        x"6400",
        x"7369",
        x"6600",
        x"756C",
        x"6873",
        x"6600",
        x"6C69",
        x"006C",
        x"7263",
        x"0063",
        x"6F63",
        x"7970",
        x"6300",
        x"6D6F",
        x"6170",
        x"6572",
        x"6D00",
        x"6D65",
        x"7700",
        x"0072",
        x"6F67",
        x"6500",
        x"6578",
        x"0063",
        x"6F6D",
        x"6564",
        x"7400",
        x"7365",
        x"0074",
        x"6F6C",
        x"6461",
        x"7300",
        x"7661",
        x"0065",
        x"7273",
        x"6365",
        x"7300",
        x"6570",
        x"6963",
        x"6C61",
        x"7200",
        x"7365",
        x"7465",
        x"7400",
        x"6172",
        x"6563",
        x"6200",
        x"696C",
        x"7473",
        x"6200",
        x"6572",
        x"6B61",
        x"0078",
        x"6177",
        x"6374",
        x"7868",
        x"6200",
        x"6572",
        x"6B61",
        x"0072",
        x"6177",
        x"6374",
        x"7268",
        x"6200",
        x"6572",
        x"6B61",
        x"0077",
        x"6177",
        x"6374",
        x"7768",
        x"6300",
        x"656C",
        x"7261",
        x"7400",
        x"6972",
        x"6767",
        x"7265",
        x"1B00",
        x"325B",
        x"004A",
        x"5B1B",
        x"3B30",
        x"4830",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000",
        x"0000"
    );

begin

    process (cp2)
    begin
        if rising_edge(cp2) then
            if ce = '1' then
                if (we = '1') then
                    RAM(conv_integer(address)) <= din;
                end if;
                dout <= RAM(conv_integer(address));
            end if;
        end if;
    end process;

end RTL;
